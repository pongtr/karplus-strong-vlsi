magic
tech scmos
timestamp 1037203521
<< ndiffusion >>
rect 12 98 17 102
rect 21 98 27 102
rect 31 98 37 102
rect 41 98 47 102
rect 51 98 56 102
rect 12 97 56 98
rect 16 93 22 97
rect 26 93 32 97
rect 36 93 42 97
rect 46 93 52 97
rect 12 92 56 93
rect 12 88 17 92
rect 21 88 27 92
rect 31 88 37 92
rect 41 88 47 92
rect 51 88 56 92
rect 12 87 56 88
rect 16 83 22 87
rect 26 83 32 87
rect 36 83 42 87
rect 46 83 52 87
rect 12 82 56 83
rect 12 78 17 82
rect 21 78 27 82
rect 31 78 37 82
rect 41 78 47 82
rect 51 78 56 82
rect 12 77 56 78
rect 16 73 22 77
rect 26 73 32 77
rect 36 73 42 77
rect 46 73 52 77
rect 12 72 56 73
rect 12 68 17 72
rect 21 68 27 72
rect 31 68 37 72
rect 41 68 47 72
rect 51 68 56 72
rect 12 67 56 68
rect 16 63 22 67
rect 26 63 32 67
rect 36 63 42 67
rect 46 63 52 67
rect 12 62 56 63
rect 12 58 17 62
rect 21 58 27 62
rect 31 58 37 62
rect 41 58 47 62
rect 51 58 56 62
rect 12 57 56 58
rect 16 53 22 57
rect 26 53 32 57
rect 36 53 42 57
rect 46 53 52 57
rect 12 52 56 53
rect 12 48 17 52
rect 21 48 27 52
rect 31 48 37 52
rect 41 48 47 52
rect 51 48 56 52
rect 12 47 56 48
rect 16 43 22 47
rect 26 43 32 47
rect 36 43 42 47
rect 46 43 52 47
rect 12 42 56 43
rect 12 38 17 42
rect 21 38 27 42
rect 31 38 37 42
rect 41 38 47 42
rect 51 38 56 42
rect 12 37 56 38
rect 16 33 22 37
rect 26 33 32 37
rect 36 33 42 37
rect 46 33 52 37
rect 12 32 56 33
rect 12 28 17 32
rect 21 28 27 32
rect 31 28 37 32
rect 41 28 47 32
rect 51 28 56 32
rect 12 27 56 28
rect 16 23 22 27
rect 26 23 32 27
rect 36 23 42 27
rect 46 23 52 27
rect 12 22 56 23
rect 12 18 17 22
rect 21 18 27 22
rect 31 18 37 22
rect 41 18 47 22
rect 51 18 56 22
rect 12 17 56 18
rect 16 13 22 17
rect 26 13 32 17
rect 36 13 42 17
rect 46 13 52 17
<< ndcontact >>
rect 17 98 21 102
rect 27 98 31 102
rect 37 98 41 102
rect 47 98 51 102
rect 12 93 16 97
rect 22 93 26 97
rect 32 93 36 97
rect 42 93 46 97
rect 52 93 56 97
rect 17 88 21 92
rect 27 88 31 92
rect 37 88 41 92
rect 47 88 51 92
rect 12 83 16 87
rect 22 83 26 87
rect 32 83 36 87
rect 42 83 46 87
rect 52 83 56 87
rect 17 78 21 82
rect 27 78 31 82
rect 37 78 41 82
rect 47 78 51 82
rect 12 73 16 77
rect 22 73 26 77
rect 32 73 36 77
rect 42 73 46 77
rect 52 73 56 77
rect 17 68 21 72
rect 27 68 31 72
rect 37 68 41 72
rect 47 68 51 72
rect 12 63 16 67
rect 22 63 26 67
rect 32 63 36 67
rect 42 63 46 67
rect 52 63 56 67
rect 17 58 21 62
rect 27 58 31 62
rect 37 58 41 62
rect 47 58 51 62
rect 12 53 16 57
rect 22 53 26 57
rect 32 53 36 57
rect 42 53 46 57
rect 52 53 56 57
rect 17 48 21 52
rect 27 48 31 52
rect 37 48 41 52
rect 47 48 51 52
rect 12 43 16 47
rect 22 43 26 47
rect 32 43 36 47
rect 42 43 46 47
rect 52 43 56 47
rect 17 38 21 42
rect 27 38 31 42
rect 37 38 41 42
rect 47 38 51 42
rect 12 33 16 37
rect 22 33 26 37
rect 32 33 36 37
rect 42 33 46 37
rect 52 33 56 37
rect 17 28 21 32
rect 27 28 31 32
rect 37 28 41 32
rect 47 28 51 32
rect 12 23 16 27
rect 22 23 26 27
rect 32 23 36 27
rect 42 23 46 27
rect 52 23 56 27
rect 17 18 21 22
rect 27 18 31 22
rect 37 18 41 22
rect 47 18 51 22
rect 12 13 16 17
rect 22 13 26 17
rect 32 13 36 17
rect 42 13 46 17
rect 52 13 56 17
<< psubstratepdiff >>
rect -2 114 70 116
rect -2 110 0 114
rect 4 110 7 114
rect 11 110 12 114
rect 16 110 17 114
rect 21 110 22 114
rect 26 110 27 114
rect 31 110 32 114
rect 36 110 37 114
rect 41 110 42 114
rect 46 110 47 114
rect 51 110 52 114
rect 56 110 57 114
rect 61 110 64 114
rect 68 110 70 114
rect -2 108 70 110
rect -2 107 6 108
rect -2 103 0 107
rect 4 103 6 107
rect -2 102 6 103
rect 62 107 70 108
rect 62 103 64 107
rect 68 103 70 107
rect 62 102 70 103
rect -2 98 0 102
rect 4 98 6 102
rect -2 97 6 98
rect -2 93 0 97
rect 4 93 6 97
rect -2 92 6 93
rect -2 88 0 92
rect 4 88 6 92
rect -2 87 6 88
rect -2 83 0 87
rect 4 83 6 87
rect -2 82 6 83
rect -2 78 0 82
rect 4 78 6 82
rect -2 77 6 78
rect -2 73 0 77
rect 4 73 6 77
rect -2 72 6 73
rect -2 68 0 72
rect 4 68 6 72
rect -2 67 6 68
rect -2 63 0 67
rect 4 63 6 67
rect -2 62 6 63
rect -2 58 0 62
rect 4 58 6 62
rect -2 57 6 58
rect -2 53 0 57
rect 4 53 6 57
rect -2 52 6 53
rect -2 48 0 52
rect 4 48 6 52
rect -2 47 6 48
rect -2 43 0 47
rect 4 43 6 47
rect -2 42 6 43
rect -2 38 0 42
rect 4 38 6 42
rect -2 37 6 38
rect -2 33 0 37
rect 4 33 6 37
rect -2 32 6 33
rect -2 28 0 32
rect 4 28 6 32
rect -2 27 6 28
rect -2 23 0 27
rect 4 23 6 27
rect -2 22 6 23
rect -2 18 0 22
rect 4 18 6 22
rect -2 17 6 18
rect -2 13 0 17
rect 4 13 6 17
rect 62 98 64 102
rect 68 98 70 102
rect 62 97 70 98
rect 62 93 64 97
rect 68 93 70 97
rect 62 92 70 93
rect 62 88 64 92
rect 68 88 70 92
rect 62 87 70 88
rect 62 83 64 87
rect 68 83 70 87
rect 62 82 70 83
rect 62 78 64 82
rect 68 78 70 82
rect 62 77 70 78
rect 62 73 64 77
rect 68 73 70 77
rect 62 72 70 73
rect 62 68 64 72
rect 68 68 70 72
rect 62 67 70 68
rect 62 63 64 67
rect 68 63 70 67
rect 62 62 70 63
rect 62 58 64 62
rect 68 58 70 62
rect 62 57 70 58
rect 62 53 64 57
rect 68 53 70 57
rect 62 52 70 53
rect 62 48 64 52
rect 68 48 70 52
rect 62 47 70 48
rect 62 43 64 47
rect 68 43 70 47
rect 62 42 70 43
rect 62 38 64 42
rect 68 38 70 42
rect 62 37 70 38
rect 62 33 64 37
rect 68 33 70 37
rect 62 32 70 33
rect 62 28 64 32
rect 68 28 70 32
rect 62 27 70 28
rect 62 23 64 27
rect 68 23 70 27
rect 62 22 70 23
rect 62 18 64 22
rect 68 18 70 22
rect 62 17 70 18
rect 62 13 64 17
rect 68 13 70 17
rect -2 12 6 13
rect -2 8 0 12
rect 4 8 6 12
rect -2 7 6 8
rect 62 12 70 13
rect 62 8 64 12
rect 68 8 70 12
rect 62 7 70 8
rect -2 5 70 7
rect -2 1 0 5
rect 4 1 7 5
rect 11 1 12 5
rect 16 1 17 5
rect 21 1 22 5
rect 26 1 27 5
rect 31 1 32 5
rect 36 1 37 5
rect 41 1 42 5
rect 46 1 47 5
rect 51 1 52 5
rect 56 1 57 5
rect 61 1 64 5
rect 68 1 70 5
rect -2 -1 70 1
<< nsubstratendiff >>
rect -14 127 82 128
rect -14 123 -13 127
rect -9 123 -8 127
rect -4 123 -3 127
rect 1 123 2 127
rect 6 123 7 127
rect 11 123 12 127
rect 16 123 17 127
rect 21 123 22 127
rect 26 123 27 127
rect 31 123 32 127
rect 36 123 37 127
rect 41 123 42 127
rect 46 123 47 127
rect 51 123 52 127
rect 56 123 57 127
rect 61 123 62 127
rect 66 123 67 127
rect 71 123 72 127
rect 76 123 77 127
rect 81 123 82 127
rect -14 122 82 123
rect -14 118 -13 122
rect -9 118 -8 122
rect -14 117 -8 118
rect -14 113 -13 117
rect -9 113 -8 117
rect 76 118 77 122
rect 81 118 82 122
rect 76 117 82 118
rect -14 112 -8 113
rect -14 108 -13 112
rect -9 108 -8 112
rect -14 107 -8 108
rect -14 103 -13 107
rect -9 103 -8 107
rect -14 102 -8 103
rect -14 98 -13 102
rect -9 98 -8 102
rect -14 97 -8 98
rect -14 93 -13 97
rect -9 93 -8 97
rect -14 92 -8 93
rect -14 88 -13 92
rect -9 88 -8 92
rect -14 87 -8 88
rect -14 83 -13 87
rect -9 83 -8 87
rect -14 82 -8 83
rect -14 78 -13 82
rect -9 78 -8 82
rect -14 77 -8 78
rect -14 73 -13 77
rect -9 73 -8 77
rect -14 72 -8 73
rect -14 68 -13 72
rect -9 68 -8 72
rect -14 67 -8 68
rect -14 63 -13 67
rect -9 63 -8 67
rect -14 62 -8 63
rect -14 58 -13 62
rect -9 58 -8 62
rect -14 57 -8 58
rect -14 53 -13 57
rect -9 53 -8 57
rect -14 52 -8 53
rect -14 48 -13 52
rect -9 48 -8 52
rect -14 47 -8 48
rect -14 43 -13 47
rect -9 43 -8 47
rect -14 42 -8 43
rect -14 38 -13 42
rect -9 38 -8 42
rect -14 37 -8 38
rect -14 33 -13 37
rect -9 33 -8 37
rect -14 32 -8 33
rect -14 28 -13 32
rect -9 28 -8 32
rect -14 27 -8 28
rect -14 23 -13 27
rect -9 23 -8 27
rect -14 22 -8 23
rect -14 18 -13 22
rect -9 18 -8 22
rect -14 17 -8 18
rect -14 13 -13 17
rect -9 13 -8 17
rect -14 12 -8 13
rect -14 8 -13 12
rect -9 8 -8 12
rect -14 7 -8 8
rect -14 3 -13 7
rect -9 3 -8 7
rect -14 2 -8 3
rect -14 -2 -13 2
rect -9 -2 -8 2
rect 76 113 77 117
rect 81 113 82 117
rect 76 112 82 113
rect 76 108 77 112
rect 81 108 82 112
rect 76 107 82 108
rect 76 103 77 107
rect 81 103 82 107
rect 76 102 82 103
rect 76 98 77 102
rect 81 98 82 102
rect 76 97 82 98
rect 76 93 77 97
rect 81 93 82 97
rect 76 92 82 93
rect 76 88 77 92
rect 81 88 82 92
rect 76 87 82 88
rect 76 83 77 87
rect 81 83 82 87
rect 76 82 82 83
rect 76 78 77 82
rect 81 78 82 82
rect 76 77 82 78
rect 76 73 77 77
rect 81 73 82 77
rect 76 72 82 73
rect 76 68 77 72
rect 81 68 82 72
rect 76 67 82 68
rect 76 63 77 67
rect 81 63 82 67
rect 76 62 82 63
rect 76 58 77 62
rect 81 58 82 62
rect 76 57 82 58
rect 76 53 77 57
rect 81 53 82 57
rect 76 52 82 53
rect 76 48 77 52
rect 81 48 82 52
rect 76 47 82 48
rect 76 43 77 47
rect 81 43 82 47
rect 76 42 82 43
rect 76 38 77 42
rect 81 38 82 42
rect 76 37 82 38
rect 76 33 77 37
rect 81 33 82 37
rect 76 32 82 33
rect 76 28 77 32
rect 81 28 82 32
rect 76 27 82 28
rect 76 23 77 27
rect 81 23 82 27
rect 76 22 82 23
rect 76 18 77 22
rect 81 18 82 22
rect 76 17 82 18
rect 76 13 77 17
rect 81 13 82 17
rect 76 12 82 13
rect 76 8 77 12
rect 81 8 82 12
rect 76 7 82 8
rect 76 3 77 7
rect 81 3 82 7
rect 76 2 82 3
rect -14 -3 -8 -2
rect -14 -7 -13 -3
rect -9 -7 -8 -3
rect 76 -2 77 2
rect 81 -2 82 2
rect 76 -3 82 -2
rect 76 -7 77 -3
rect 81 -7 82 -3
rect -14 -8 82 -7
rect -14 -12 -13 -8
rect -9 -12 -8 -8
rect -4 -12 -3 -8
rect 1 -12 2 -8
rect 6 -12 7 -8
rect 11 -12 12 -8
rect 16 -12 17 -8
rect 21 -12 22 -8
rect 26 -12 27 -8
rect 31 -12 32 -8
rect 36 -12 37 -8
rect 41 -12 42 -8
rect 46 -12 47 -8
rect 51 -12 52 -8
rect 56 -12 57 -8
rect 61 -12 62 -8
rect 66 -12 67 -8
rect 71 -12 72 -8
rect 76 -12 77 -8
rect 81 -12 82 -8
rect -14 -13 82 -12
<< psubstratepcontact >>
rect 0 110 4 114
rect 7 110 11 114
rect 12 110 16 114
rect 17 110 21 114
rect 22 110 26 114
rect 27 110 31 114
rect 32 110 36 114
rect 37 110 41 114
rect 42 110 46 114
rect 47 110 51 114
rect 52 110 56 114
rect 57 110 61 114
rect 64 110 68 114
rect 0 103 4 107
rect 64 103 68 107
rect 0 98 4 102
rect 0 93 4 97
rect 0 88 4 92
rect 0 83 4 87
rect 0 78 4 82
rect 0 73 4 77
rect 0 68 4 72
rect 0 63 4 67
rect 0 58 4 62
rect 0 53 4 57
rect 0 48 4 52
rect 0 43 4 47
rect 0 38 4 42
rect 0 33 4 37
rect 0 28 4 32
rect 0 23 4 27
rect 0 18 4 22
rect 0 13 4 17
rect 64 98 68 102
rect 64 93 68 97
rect 64 88 68 92
rect 64 83 68 87
rect 64 78 68 82
rect 64 73 68 77
rect 64 68 68 72
rect 64 63 68 67
rect 64 58 68 62
rect 64 53 68 57
rect 64 48 68 52
rect 64 43 68 47
rect 64 38 68 42
rect 64 33 68 37
rect 64 28 68 32
rect 64 23 68 27
rect 64 18 68 22
rect 64 13 68 17
rect 0 8 4 12
rect 64 8 68 12
rect 0 1 4 5
rect 7 1 11 5
rect 12 1 16 5
rect 17 1 21 5
rect 22 1 26 5
rect 27 1 31 5
rect 32 1 36 5
rect 37 1 41 5
rect 42 1 46 5
rect 47 1 51 5
rect 52 1 56 5
rect 57 1 61 5
rect 64 1 68 5
<< nsubstratencontact >>
rect -13 123 -9 127
rect -8 123 -4 127
rect -3 123 1 127
rect 2 123 6 127
rect 7 123 11 127
rect 12 123 16 127
rect 17 123 21 127
rect 22 123 26 127
rect 27 123 31 127
rect 32 123 36 127
rect 37 123 41 127
rect 42 123 46 127
rect 47 123 51 127
rect 52 123 56 127
rect 57 123 61 127
rect 62 123 66 127
rect 67 123 71 127
rect 72 123 76 127
rect 77 123 81 127
rect -13 118 -9 122
rect -13 113 -9 117
rect 77 118 81 122
rect -13 108 -9 112
rect -13 103 -9 107
rect -13 98 -9 102
rect -13 93 -9 97
rect -13 88 -9 92
rect -13 83 -9 87
rect -13 78 -9 82
rect -13 73 -9 77
rect -13 68 -9 72
rect -13 63 -9 67
rect -13 58 -9 62
rect -13 53 -9 57
rect -13 48 -9 52
rect -13 43 -9 47
rect -13 38 -9 42
rect -13 33 -9 37
rect -13 28 -9 32
rect -13 23 -9 27
rect -13 18 -9 22
rect -13 13 -9 17
rect -13 8 -9 12
rect -13 3 -9 7
rect -13 -2 -9 2
rect 77 113 81 117
rect 77 108 81 112
rect 77 103 81 107
rect 77 98 81 102
rect 77 93 81 97
rect 77 88 81 92
rect 77 83 81 87
rect 77 78 81 82
rect 77 73 81 77
rect 77 68 81 72
rect 77 63 81 67
rect 77 58 81 62
rect 77 53 81 57
rect 77 48 81 52
rect 77 43 81 47
rect 77 38 81 42
rect 77 33 81 37
rect 77 28 81 32
rect 77 23 81 27
rect 77 18 81 22
rect 77 13 81 17
rect 77 8 81 12
rect 77 3 81 7
rect -13 -7 -9 -3
rect 77 -2 81 2
rect 77 -7 81 -3
rect -13 -12 -9 -8
rect -8 -12 -4 -8
rect -3 -12 1 -8
rect 2 -12 6 -8
rect 7 -12 11 -8
rect 12 -12 16 -8
rect 17 -12 21 -8
rect 22 -12 26 -8
rect 27 -12 31 -8
rect 32 -12 36 -8
rect 37 -12 41 -8
rect 42 -12 46 -8
rect 47 -12 51 -8
rect 52 -12 56 -8
rect 57 -12 61 -8
rect 62 -12 66 -8
rect 67 -12 71 -8
rect 72 -12 76 -8
rect 77 -12 81 -8
<< metal1 >>
rect -9 123 -8 127
rect -4 123 -3 127
rect 1 123 2 127
rect 6 123 7 127
rect 11 123 12 127
rect 16 123 17 127
rect 21 123 22 127
rect 26 123 27 127
rect 31 123 32 127
rect 36 123 37 127
rect 41 123 42 127
rect 46 123 47 127
rect 51 123 52 127
rect 56 123 57 127
rect 61 123 62 127
rect 66 123 67 127
rect 71 123 72 127
rect 76 123 77 127
rect -13 122 -9 123
rect -13 117 -9 118
rect 77 122 81 123
rect 77 117 81 118
rect -13 112 -9 113
rect -13 107 -9 108
rect -13 102 -9 103
rect -13 97 -9 98
rect -13 92 -9 93
rect -13 87 -9 88
rect -13 82 -9 83
rect -13 77 -9 78
rect -13 72 -9 73
rect -13 67 -9 68
rect -13 62 -9 63
rect -13 57 -9 58
rect -13 52 -9 53
rect -13 47 -9 48
rect -13 42 -9 43
rect -13 37 -9 38
rect -13 32 -9 33
rect -13 27 -9 28
rect -13 22 -9 23
rect -13 17 -9 18
rect -13 12 -9 13
rect -13 7 -9 8
rect -13 2 -9 3
rect 4 110 7 114
rect 11 110 12 114
rect 16 110 17 114
rect 21 110 22 114
rect 26 110 27 114
rect 31 110 32 114
rect 36 110 37 114
rect 41 110 42 114
rect 46 110 47 114
rect 51 110 52 114
rect 56 110 57 114
rect 61 110 64 114
rect 0 107 4 110
rect 0 102 4 103
rect 64 107 68 110
rect 64 102 68 103
rect 0 97 4 98
rect 0 92 4 93
rect 0 87 4 88
rect 0 82 4 83
rect 0 77 4 78
rect 0 72 4 73
rect 0 67 4 68
rect 0 62 4 63
rect 0 57 4 58
rect 0 52 4 53
rect 0 47 4 48
rect 0 42 4 43
rect 0 37 4 38
rect 0 32 4 33
rect 0 27 4 28
rect 0 22 4 23
rect 0 17 4 18
rect 16 98 17 102
rect 21 98 22 102
rect 26 98 27 102
rect 31 98 32 102
rect 36 98 37 102
rect 41 98 42 102
rect 46 98 47 102
rect 51 98 52 102
rect 12 97 56 98
rect 16 93 17 97
rect 21 93 22 97
rect 26 93 27 97
rect 31 93 32 97
rect 36 93 37 97
rect 41 93 42 97
rect 46 93 47 97
rect 51 93 52 97
rect 12 92 56 93
rect 16 88 17 92
rect 21 88 22 92
rect 26 88 27 92
rect 31 88 32 92
rect 36 88 37 92
rect 41 88 42 92
rect 46 88 47 92
rect 51 88 52 92
rect 12 87 56 88
rect 16 83 17 87
rect 21 83 22 87
rect 26 83 27 87
rect 31 83 32 87
rect 36 83 37 87
rect 41 83 42 87
rect 46 83 47 87
rect 51 83 52 87
rect 12 82 56 83
rect 16 78 17 82
rect 21 78 22 82
rect 26 78 27 82
rect 31 78 32 82
rect 36 78 37 82
rect 41 78 42 82
rect 46 78 47 82
rect 51 78 52 82
rect 12 77 56 78
rect 16 73 17 77
rect 21 73 22 77
rect 26 73 27 77
rect 31 73 32 77
rect 36 73 37 77
rect 41 73 42 77
rect 46 73 47 77
rect 51 73 52 77
rect 12 72 56 73
rect 16 68 17 72
rect 21 68 22 72
rect 26 68 27 72
rect 31 68 32 72
rect 36 68 37 72
rect 41 68 42 72
rect 46 68 47 72
rect 51 68 52 72
rect 12 67 56 68
rect 16 63 17 67
rect 21 63 22 67
rect 26 63 27 67
rect 31 63 32 67
rect 36 63 37 67
rect 41 63 42 67
rect 46 63 47 67
rect 51 63 52 67
rect 12 62 56 63
rect 16 58 17 62
rect 21 58 22 62
rect 26 58 27 62
rect 31 58 32 62
rect 36 58 37 62
rect 41 58 42 62
rect 46 58 47 62
rect 51 58 52 62
rect 12 57 56 58
rect 16 53 17 57
rect 21 53 22 57
rect 26 53 27 57
rect 31 53 32 57
rect 36 53 37 57
rect 41 53 42 57
rect 46 53 47 57
rect 51 53 52 57
rect 12 52 56 53
rect 16 48 17 52
rect 21 48 22 52
rect 26 48 27 52
rect 31 48 32 52
rect 36 48 37 52
rect 41 48 42 52
rect 46 48 47 52
rect 51 48 52 52
rect 12 47 56 48
rect 16 43 17 47
rect 21 43 22 47
rect 26 43 27 47
rect 31 43 32 47
rect 36 43 37 47
rect 41 43 42 47
rect 46 43 47 47
rect 51 43 52 47
rect 12 42 56 43
rect 16 38 17 42
rect 21 38 22 42
rect 26 38 27 42
rect 31 38 32 42
rect 36 38 37 42
rect 41 38 42 42
rect 46 38 47 42
rect 51 38 52 42
rect 12 37 56 38
rect 16 33 17 37
rect 21 33 22 37
rect 26 33 27 37
rect 31 33 32 37
rect 36 33 37 37
rect 41 33 42 37
rect 46 33 47 37
rect 51 33 52 37
rect 12 32 56 33
rect 16 28 17 32
rect 21 28 22 32
rect 26 28 27 32
rect 31 28 32 32
rect 36 28 37 32
rect 41 28 42 32
rect 46 28 47 32
rect 51 28 52 32
rect 12 27 56 28
rect 16 23 17 27
rect 21 23 22 27
rect 26 23 27 27
rect 31 23 32 27
rect 36 23 37 27
rect 41 23 42 27
rect 46 23 47 27
rect 51 23 52 27
rect 12 22 56 23
rect 16 18 17 22
rect 21 18 22 22
rect 26 18 27 22
rect 31 18 32 22
rect 36 18 37 22
rect 41 18 42 22
rect 46 18 47 22
rect 51 18 52 22
rect 12 17 56 18
rect 16 13 17 17
rect 21 13 22 17
rect 26 13 27 17
rect 31 13 32 17
rect 36 13 37 17
rect 41 13 42 17
rect 46 13 47 17
rect 51 13 52 17
rect 64 97 68 98
rect 64 92 68 93
rect 64 87 68 88
rect 64 82 68 83
rect 64 77 68 78
rect 64 72 68 73
rect 64 67 68 68
rect 64 62 68 63
rect 64 57 68 58
rect 64 52 68 53
rect 64 47 68 48
rect 64 42 68 43
rect 64 37 68 38
rect 64 32 68 33
rect 64 27 68 28
rect 64 22 68 23
rect 64 17 68 18
rect 0 12 4 13
rect 0 5 4 8
rect 64 12 68 13
rect 64 5 68 8
rect 4 1 7 5
rect 11 1 12 5
rect 16 1 17 5
rect 21 1 22 5
rect 26 1 27 5
rect 31 1 32 5
rect 36 1 37 5
rect 41 1 42 5
rect 46 1 47 5
rect 51 1 52 5
rect 56 1 57 5
rect 61 1 64 5
rect 77 112 81 113
rect 77 107 81 108
rect 77 102 81 103
rect 77 97 81 98
rect 77 92 81 93
rect 77 87 81 88
rect 77 82 81 83
rect 77 77 81 78
rect 77 72 81 73
rect 77 67 81 68
rect 77 62 81 63
rect 77 57 81 58
rect 77 52 81 53
rect 77 47 81 48
rect 77 42 81 43
rect 77 37 81 38
rect 77 32 81 33
rect 77 27 81 28
rect 77 22 81 23
rect 77 17 81 18
rect 77 12 81 13
rect 77 7 81 8
rect 77 2 81 3
rect -13 -3 -9 -2
rect -13 -8 -9 -7
rect 77 -3 81 -2
rect 77 -8 81 -7
rect -9 -12 -8 -8
rect -4 -12 -3 -8
rect 1 -12 2 -8
rect 6 -12 7 -8
rect 11 -12 12 -8
rect 16 -12 17 -8
rect 21 -12 22 -8
rect 26 -12 27 -8
rect 31 -12 32 -8
rect 36 -12 37 -8
rect 41 -12 42 -8
rect 46 -12 47 -8
rect 51 -12 52 -8
rect 56 -12 57 -8
rect 61 -12 62 -8
rect 66 -12 67 -8
rect 71 -12 72 -8
rect 76 -12 77 -8
<< m2contact >>
rect 12 98 16 102
rect 22 98 26 102
rect 32 98 36 102
rect 42 98 46 102
rect 52 98 56 102
rect 17 93 21 97
rect 27 93 31 97
rect 37 93 41 97
rect 47 93 51 97
rect 12 88 16 92
rect 22 88 26 92
rect 32 88 36 92
rect 42 88 46 92
rect 52 88 56 92
rect 17 83 21 87
rect 27 83 31 87
rect 37 83 41 87
rect 47 83 51 87
rect 12 78 16 82
rect 22 78 26 82
rect 32 78 36 82
rect 42 78 46 82
rect 52 78 56 82
rect 17 73 21 77
rect 27 73 31 77
rect 37 73 41 77
rect 47 73 51 77
rect 12 68 16 72
rect 22 68 26 72
rect 32 68 36 72
rect 42 68 46 72
rect 52 68 56 72
rect 17 63 21 67
rect 27 63 31 67
rect 37 63 41 67
rect 47 63 51 67
rect 12 58 16 62
rect 22 58 26 62
rect 32 58 36 62
rect 42 58 46 62
rect 52 58 56 62
rect 17 53 21 57
rect 27 53 31 57
rect 37 53 41 57
rect 47 53 51 57
rect 12 48 16 52
rect 22 48 26 52
rect 32 48 36 52
rect 42 48 46 52
rect 52 48 56 52
rect 17 43 21 47
rect 27 43 31 47
rect 37 43 41 47
rect 47 43 51 47
rect 12 38 16 42
rect 22 38 26 42
rect 32 38 36 42
rect 42 38 46 42
rect 52 38 56 42
rect 17 33 21 37
rect 27 33 31 37
rect 37 33 41 37
rect 47 33 51 37
rect 12 28 16 32
rect 22 28 26 32
rect 32 28 36 32
rect 42 28 46 32
rect 52 28 56 32
rect 17 23 21 27
rect 27 23 31 27
rect 37 23 41 27
rect 47 23 51 27
rect 12 18 16 22
rect 22 18 26 22
rect 32 18 36 22
rect 42 18 46 22
rect 52 18 56 22
rect 17 13 21 17
rect 27 13 31 17
rect 37 13 41 17
rect 47 13 51 17
<< metal2 >>
rect 16 98 22 102
rect 26 98 32 102
rect 36 98 42 102
rect 46 98 52 102
rect 12 97 56 98
rect 12 93 17 97
rect 21 93 27 97
rect 31 93 37 97
rect 41 93 47 97
rect 51 93 56 97
rect 12 92 56 93
rect 16 88 22 92
rect 26 88 32 92
rect 36 88 42 92
rect 46 88 52 92
rect 12 87 56 88
rect 12 83 17 87
rect 21 83 27 87
rect 31 83 37 87
rect 41 83 47 87
rect 51 83 56 87
rect 12 82 56 83
rect 16 78 22 82
rect 26 78 32 82
rect 36 78 42 82
rect 46 78 52 82
rect 12 77 56 78
rect 12 73 17 77
rect 21 73 27 77
rect 31 73 37 77
rect 41 73 47 77
rect 51 73 56 77
rect 12 72 56 73
rect 16 68 22 72
rect 26 68 32 72
rect 36 68 42 72
rect 46 68 52 72
rect 12 67 56 68
rect 12 63 17 67
rect 21 63 27 67
rect 31 63 37 67
rect 41 63 47 67
rect 51 63 56 67
rect 12 62 56 63
rect 16 58 22 62
rect 26 58 32 62
rect 36 58 42 62
rect 46 58 52 62
rect 12 57 56 58
rect 12 53 17 57
rect 21 53 27 57
rect 31 53 37 57
rect 41 53 47 57
rect 51 53 56 57
rect 12 52 56 53
rect 16 48 22 52
rect 26 48 32 52
rect 36 48 42 52
rect 46 48 52 52
rect 12 47 56 48
rect 12 43 17 47
rect 21 43 27 47
rect 31 43 37 47
rect 41 43 47 47
rect 51 43 56 47
rect 12 42 56 43
rect 16 38 22 42
rect 26 38 32 42
rect 36 38 42 42
rect 46 38 52 42
rect 12 37 56 38
rect 12 33 17 37
rect 21 33 27 37
rect 31 33 37 37
rect 41 33 47 37
rect 51 33 56 37
rect 12 32 56 33
rect 16 28 22 32
rect 26 28 32 32
rect 36 28 42 32
rect 46 28 52 32
rect 12 27 56 28
rect 12 23 17 27
rect 21 23 27 27
rect 31 23 37 27
rect 41 23 47 27
rect 51 23 56 27
rect 12 22 56 23
rect 16 18 22 22
rect 26 18 32 22
rect 36 18 42 22
rect 46 18 52 22
rect 12 17 56 18
rect 12 13 17 17
rect 21 13 27 17
rect 31 13 37 17
rect 41 13 47 17
rect 51 13 56 17
<< end >>
