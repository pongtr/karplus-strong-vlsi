magic
tech scmos
timestamp 1509371954
<< nsubstratendiff >>
rect 144 94 150 125
rect 159 94 165 125
<< metal1 >>
rect 97 356 213 357
rect 97 352 110 356
rect 114 352 117 356
rect 121 352 124 356
rect 128 352 131 356
rect 135 352 138 356
rect 142 352 145 356
rect 149 352 152 356
rect 156 352 159 356
rect 163 352 166 356
rect 170 352 173 356
rect 177 352 180 356
rect 184 352 187 356
rect 191 352 194 356
rect 198 352 213 356
rect 97 351 213 352
rect 97 348 110 351
rect 107 347 110 348
rect 114 347 117 351
rect 121 347 124 351
rect 128 347 131 351
rect 135 347 138 351
rect 142 347 145 351
rect 149 347 152 351
rect 156 347 159 351
rect 163 347 166 351
rect 170 347 173 351
rect 177 347 180 351
rect 184 347 187 351
rect 191 347 194 351
rect 198 348 213 351
rect 198 347 203 348
rect 107 346 203 347
rect 107 342 110 346
rect 114 342 117 346
rect 121 342 124 346
rect 128 342 131 346
rect 135 342 138 346
rect 142 342 145 346
rect 149 342 152 346
rect 156 342 159 346
rect 163 342 166 346
rect 170 342 173 346
rect 177 342 180 346
rect 184 342 187 346
rect 191 342 194 346
rect 198 342 203 346
rect 107 341 203 342
rect 107 337 110 341
rect 114 337 117 341
rect 121 337 124 341
rect 128 337 131 341
rect 135 337 138 341
rect 142 337 145 341
rect 149 337 152 341
rect 156 337 159 341
rect 163 337 166 341
rect 170 337 173 341
rect 177 337 180 341
rect 184 337 187 341
rect 191 337 194 341
rect 198 337 203 341
rect 107 336 203 337
rect 45 203 48 207
rect 52 203 53 207
rect 57 203 58 207
rect 62 203 63 207
rect 67 203 68 207
rect 72 203 73 207
rect 77 203 78 207
rect 82 203 83 207
rect 87 203 88 207
rect 92 203 93 207
rect 97 203 98 207
rect 102 203 105 207
rect 31 157 87 194
rect 19 155 87 157
rect 19 151 20 155
rect 24 151 25 155
rect 29 151 87 155
rect 19 150 87 151
rect 19 146 20 150
rect 24 146 25 150
rect 29 146 87 150
rect 19 145 87 146
rect 19 141 20 145
rect 24 141 25 145
rect 29 141 87 145
rect 19 140 87 141
rect 19 136 20 140
rect 24 136 25 140
rect 29 136 87 140
rect 19 135 87 136
rect 19 131 20 135
rect 24 131 25 135
rect 29 131 87 135
rect 19 130 87 131
rect 19 126 20 130
rect 24 126 25 130
rect 29 126 87 130
rect 19 125 87 126
rect 19 121 20 125
rect 24 121 25 125
rect 29 121 87 125
rect 19 120 87 121
rect 19 116 20 120
rect 24 116 25 120
rect 29 116 87 120
rect 19 115 87 116
rect 19 111 20 115
rect 24 111 25 115
rect 29 111 87 115
rect 19 110 87 111
rect 19 106 20 110
rect 24 106 25 110
rect 29 106 87 110
rect 19 105 87 106
rect 19 101 20 105
rect 24 101 25 105
rect 29 101 87 105
rect 19 100 87 101
rect 19 96 20 100
rect 24 96 25 100
rect 29 96 87 100
rect 19 95 87 96
rect 19 91 20 95
rect 24 91 25 95
rect 29 91 87 95
rect 19 89 87 91
rect 127 150 181 336
rect 205 203 208 207
rect 212 203 213 207
rect 217 203 218 207
rect 222 203 223 207
rect 227 203 228 207
rect 232 203 233 207
rect 237 203 238 207
rect 242 203 243 207
rect 247 203 248 207
rect 252 203 253 207
rect 257 203 258 207
rect 262 203 265 207
rect 127 146 155 150
rect 159 146 160 150
rect 164 146 181 150
rect 127 145 181 146
rect 127 141 155 145
rect 159 141 160 145
rect 164 141 181 145
rect 127 140 181 141
rect 127 136 155 140
rect 159 136 160 140
rect 164 136 181 140
rect 127 135 181 136
rect 127 131 155 135
rect 159 131 160 135
rect 164 131 181 135
rect 127 130 181 131
rect 127 126 155 130
rect 159 126 160 130
rect 164 126 181 130
rect 127 125 181 126
rect 127 121 155 125
rect 159 121 160 125
rect 164 121 181 125
rect 127 120 181 121
rect 127 116 155 120
rect 159 116 160 120
rect 164 116 181 120
rect 127 115 181 116
rect 127 111 155 115
rect 159 111 160 115
rect 164 111 181 115
rect 127 110 181 111
rect 127 106 155 110
rect 159 106 160 110
rect 164 106 181 110
rect 127 105 181 106
rect 127 101 155 105
rect 159 101 160 105
rect 164 101 181 105
rect 127 100 181 101
rect 127 96 155 100
rect 159 96 160 100
rect 164 96 181 100
rect 127 -35 181 96
rect 225 77 281 194
rect 229 73 230 77
rect 234 73 235 77
rect 239 73 240 77
rect 244 73 245 77
rect 249 73 250 77
rect 254 73 255 77
rect 259 73 260 77
rect 264 73 265 77
rect 269 73 270 77
rect 274 73 275 77
rect 279 73 281 77
rect 225 72 281 73
rect 229 68 230 72
rect 234 68 235 72
rect 239 68 240 72
rect 244 68 245 72
rect 249 68 250 72
rect 254 68 255 72
rect 259 68 260 72
rect 264 68 265 72
rect 269 68 270 72
rect 274 68 275 72
rect 279 68 281 72
rect 225 67 281 68
<< m2contact >>
rect 110 352 114 356
rect 117 352 121 356
rect 124 352 128 356
rect 131 352 135 356
rect 138 352 142 356
rect 145 352 149 356
rect 152 352 156 356
rect 159 352 163 356
rect 166 352 170 356
rect 173 352 177 356
rect 180 352 184 356
rect 187 352 191 356
rect 194 352 198 356
rect 110 347 114 351
rect 117 347 121 351
rect 124 347 128 351
rect 131 347 135 351
rect 138 347 142 351
rect 145 347 149 351
rect 152 347 156 351
rect 159 347 163 351
rect 166 347 170 351
rect 173 347 177 351
rect 180 347 184 351
rect 187 347 191 351
rect 194 347 198 351
rect 110 342 114 346
rect 117 342 121 346
rect 124 342 128 346
rect 131 342 135 346
rect 138 342 142 346
rect 145 342 149 346
rect 152 342 156 346
rect 159 342 163 346
rect 166 342 170 346
rect 173 342 177 346
rect 180 342 184 346
rect 187 342 191 346
rect 194 342 198 346
rect 110 337 114 341
rect 117 337 121 341
rect 124 337 128 341
rect 131 337 135 341
rect 138 337 142 341
rect 145 337 149 341
rect 152 337 156 341
rect 159 337 163 341
rect 166 337 170 341
rect 173 337 177 341
rect 180 337 184 341
rect 187 337 191 341
rect 194 337 198 341
rect 41 203 45 207
rect 48 203 52 207
rect 53 203 57 207
rect 58 203 62 207
rect 63 203 67 207
rect 68 203 72 207
rect 73 203 77 207
rect 78 203 82 207
rect 83 203 87 207
rect 88 203 92 207
rect 93 203 97 207
rect 98 203 102 207
rect 105 203 109 207
rect 20 151 24 155
rect 25 151 29 155
rect 20 146 24 150
rect 25 146 29 150
rect 20 141 24 145
rect 25 141 29 145
rect 20 136 24 140
rect 25 136 29 140
rect 20 131 24 135
rect 25 131 29 135
rect 20 126 24 130
rect 25 126 29 130
rect 20 121 24 125
rect 25 121 29 125
rect 20 116 24 120
rect 25 116 29 120
rect 20 111 24 115
rect 25 111 29 115
rect 20 106 24 110
rect 25 106 29 110
rect 20 101 24 105
rect 25 101 29 105
rect 20 96 24 100
rect 25 96 29 100
rect 20 91 24 95
rect 25 91 29 95
rect 201 203 205 207
rect 208 203 212 207
rect 213 203 217 207
rect 218 203 222 207
rect 223 203 227 207
rect 228 203 232 207
rect 233 203 237 207
rect 238 203 242 207
rect 243 203 247 207
rect 248 203 252 207
rect 253 203 257 207
rect 258 203 262 207
rect 265 203 269 207
rect 155 146 159 150
rect 160 146 164 150
rect 155 141 159 145
rect 160 141 164 145
rect 155 136 159 140
rect 160 136 164 140
rect 155 131 159 135
rect 160 131 164 135
rect 155 126 159 130
rect 160 126 164 130
rect 155 121 159 125
rect 160 121 164 125
rect 155 116 159 120
rect 160 116 164 120
rect 155 111 159 115
rect 160 111 164 115
rect 155 106 159 110
rect 160 106 164 110
rect 155 101 159 105
rect 160 101 164 105
rect 155 96 159 100
rect 160 96 164 100
rect 225 73 229 77
rect 230 73 234 77
rect 235 73 239 77
rect 240 73 244 77
rect 245 73 249 77
rect 250 73 254 77
rect 255 73 259 77
rect 260 73 264 77
rect 265 73 269 77
rect 270 73 274 77
rect 275 73 279 77
rect 225 68 229 72
rect 230 68 234 72
rect 235 68 239 72
rect 240 68 244 72
rect 245 68 249 72
rect 250 68 254 72
rect 255 68 259 72
rect 260 68 264 72
rect 265 68 269 72
rect 270 68 274 72
rect 275 68 279 72
<< metal2 >>
rect 97 356 213 357
rect 97 352 110 356
rect 114 352 117 356
rect 121 352 124 356
rect 128 352 131 356
rect 135 352 138 356
rect 142 352 145 356
rect 149 352 152 356
rect 156 352 159 356
rect 163 352 166 356
rect 170 352 173 356
rect 177 352 180 356
rect 184 352 187 356
rect 191 352 194 356
rect 198 352 213 356
rect 97 351 213 352
rect 97 348 110 351
rect 107 347 110 348
rect 114 347 117 351
rect 121 347 124 351
rect 128 347 131 351
rect 135 347 138 351
rect 142 347 145 351
rect 149 347 152 351
rect 156 347 159 351
rect 163 347 166 351
rect 170 347 173 351
rect 177 347 180 351
rect 184 347 187 351
rect 191 347 194 351
rect 198 348 213 351
rect 198 347 203 348
rect 107 346 203 347
rect 107 342 110 346
rect 114 342 117 346
rect 121 342 124 346
rect 128 342 131 346
rect 135 342 138 346
rect 142 342 145 346
rect 149 342 152 346
rect 156 342 159 346
rect 163 342 166 346
rect 170 342 173 346
rect 177 342 180 346
rect 184 342 187 346
rect 191 342 194 346
rect 198 342 203 346
rect 107 341 203 342
rect 107 337 110 341
rect 114 337 117 341
rect 121 337 124 341
rect 128 337 131 341
rect 135 337 138 341
rect 142 337 145 341
rect 149 337 152 341
rect 156 337 159 341
rect 163 337 166 341
rect 170 337 173 341
rect 177 337 180 341
rect 184 337 187 341
rect 191 337 194 341
rect 198 337 203 341
rect 107 308 203 337
rect 97 219 213 308
rect 45 203 48 207
rect 52 203 53 207
rect 57 203 58 207
rect 62 203 63 207
rect 67 203 68 207
rect 72 203 73 207
rect 77 203 78 207
rect 82 203 83 207
rect 87 203 88 207
rect 92 203 93 207
rect 97 203 98 207
rect 102 203 105 207
rect 8 155 29 157
rect 8 151 10 155
rect 14 151 15 155
rect 19 151 20 155
rect 24 151 25 155
rect 8 150 29 151
rect 8 146 10 150
rect 14 146 15 150
rect 19 146 20 150
rect 24 146 25 150
rect 8 145 29 146
rect 8 141 10 145
rect 14 141 15 145
rect 19 141 20 145
rect 24 141 25 145
rect 8 140 29 141
rect 8 136 10 140
rect 14 136 15 140
rect 19 136 20 140
rect 24 136 25 140
rect 8 135 29 136
rect 8 131 10 135
rect 14 131 15 135
rect 19 131 20 135
rect 24 131 25 135
rect 8 130 29 131
rect 8 126 10 130
rect 14 126 15 130
rect 19 126 20 130
rect 24 126 25 130
rect 8 125 29 126
rect 8 121 10 125
rect 14 121 15 125
rect 19 121 20 125
rect 24 121 25 125
rect 8 120 29 121
rect 8 116 10 120
rect 14 116 15 120
rect 19 116 20 120
rect 24 116 25 120
rect 8 115 29 116
rect 8 111 10 115
rect 14 111 15 115
rect 19 111 20 115
rect 24 111 25 115
rect 8 110 29 111
rect 8 106 10 110
rect 14 106 15 110
rect 19 106 20 110
rect 24 106 25 110
rect 8 105 29 106
rect 8 101 10 105
rect 14 101 15 105
rect 19 101 20 105
rect 24 101 25 105
rect 8 100 29 101
rect 8 96 10 100
rect 14 96 15 100
rect 19 96 20 100
rect 24 96 25 100
rect 8 95 29 96
rect 8 91 10 95
rect 14 91 15 95
rect 19 91 20 95
rect 24 91 25 95
rect 8 89 29 91
rect 41 67 109 203
rect 205 203 208 207
rect 212 203 213 207
rect 217 203 218 207
rect 222 203 223 207
rect 227 203 228 207
rect 232 203 233 207
rect 237 203 238 207
rect 242 203 243 207
rect 247 203 248 207
rect 252 203 253 207
rect 257 203 258 207
rect 262 203 265 207
rect 144 146 145 150
rect 149 146 150 150
rect 154 146 155 150
rect 159 146 160 150
rect 144 145 164 146
rect 144 141 145 145
rect 149 141 150 145
rect 154 141 155 145
rect 159 141 160 145
rect 144 140 164 141
rect 144 136 145 140
rect 149 136 150 140
rect 154 136 155 140
rect 159 136 160 140
rect 144 135 164 136
rect 144 131 145 135
rect 149 131 150 135
rect 154 131 155 135
rect 159 131 160 135
rect 144 130 164 131
rect 144 126 145 130
rect 149 126 150 130
rect 154 126 155 130
rect 159 126 160 130
rect 144 125 164 126
rect 144 121 145 125
rect 149 121 150 125
rect 154 121 155 125
rect 159 121 160 125
rect 144 120 164 121
rect 144 116 145 120
rect 149 116 150 120
rect 154 116 155 120
rect 159 116 160 120
rect 144 115 164 116
rect 144 111 145 115
rect 149 111 150 115
rect 154 111 155 115
rect 159 111 160 115
rect 201 124 269 203
rect 201 120 203 124
rect 207 120 208 124
rect 212 120 213 124
rect 217 120 218 124
rect 222 120 223 124
rect 227 120 228 124
rect 232 120 233 124
rect 237 120 238 124
rect 242 120 243 124
rect 247 120 248 124
rect 252 120 253 124
rect 257 120 258 124
rect 262 120 263 124
rect 267 120 269 124
rect 201 119 269 120
rect 201 115 203 119
rect 207 115 208 119
rect 212 115 213 119
rect 217 115 218 119
rect 222 115 223 119
rect 227 115 228 119
rect 232 115 233 119
rect 237 115 238 119
rect 242 115 243 119
rect 247 115 248 119
rect 252 115 253 119
rect 257 115 258 119
rect 262 115 263 119
rect 267 115 269 119
rect 201 112 269 115
rect 144 110 164 111
rect 144 106 145 110
rect 149 106 150 110
rect 154 106 155 110
rect 159 106 160 110
rect 144 105 164 106
rect 144 101 145 105
rect 149 101 150 105
rect 154 101 155 105
rect 159 101 160 105
rect 144 100 164 101
rect 144 96 145 100
rect 149 96 150 100
rect 154 96 155 100
rect 159 96 160 100
rect 144 94 164 96
rect 41 63 43 67
rect 47 63 48 67
rect 52 63 53 67
rect 57 63 58 67
rect 62 63 63 67
rect 67 63 68 67
rect 72 63 73 67
rect 77 63 78 67
rect 82 63 83 67
rect 87 63 88 67
rect 92 63 93 67
rect 97 63 98 67
rect 102 63 103 67
rect 107 63 109 67
rect 41 62 109 63
rect 41 58 43 62
rect 47 58 48 62
rect 52 58 53 62
rect 57 58 58 62
rect 62 58 63 62
rect 67 58 68 62
rect 72 58 73 62
rect 77 58 78 62
rect 82 58 83 62
rect 87 58 88 62
rect 92 58 93 62
rect 97 58 98 62
rect 102 58 103 62
rect 107 58 109 62
rect 41 55 109 58
rect 229 73 230 77
rect 234 73 235 77
rect 239 73 240 77
rect 244 73 245 77
rect 249 73 250 77
rect 254 73 255 77
rect 259 73 260 77
rect 264 73 265 77
rect 269 73 270 77
rect 274 73 275 77
rect 279 73 281 77
rect 225 72 281 73
rect 229 68 230 72
rect 234 68 235 72
rect 239 68 240 72
rect 244 68 245 72
rect 249 68 250 72
rect 254 68 255 72
rect 259 68 260 72
rect 264 68 265 72
rect 269 68 270 72
rect 274 68 275 72
rect 279 68 281 72
rect 225 67 281 68
rect 229 63 230 67
rect 234 63 235 67
rect 239 63 240 67
rect 244 63 245 67
rect 249 63 250 67
rect 254 63 255 67
rect 259 63 260 67
rect 264 63 265 67
rect 269 63 270 67
rect 274 63 275 67
rect 279 63 281 67
rect 225 62 281 63
rect 229 58 230 62
rect 234 58 235 62
rect 239 58 240 62
rect 244 58 245 62
rect 249 58 250 62
rect 254 58 255 62
rect 259 58 260 62
rect 264 58 265 62
rect 269 58 270 62
rect 274 58 275 62
rect 279 58 281 62
rect 225 56 281 58
<< m3contact >>
rect 10 151 14 155
rect 15 151 19 155
rect 10 146 14 150
rect 15 146 19 150
rect 10 141 14 145
rect 15 141 19 145
rect 10 136 14 140
rect 15 136 19 140
rect 10 131 14 135
rect 15 131 19 135
rect 10 126 14 130
rect 15 126 19 130
rect 10 121 14 125
rect 15 121 19 125
rect 10 116 14 120
rect 15 116 19 120
rect 10 111 14 115
rect 15 111 19 115
rect 10 106 14 110
rect 15 106 19 110
rect 10 101 14 105
rect 15 101 19 105
rect 10 96 14 100
rect 15 96 19 100
rect 10 91 14 95
rect 15 91 19 95
rect 145 146 149 150
rect 150 146 154 150
rect 145 141 149 145
rect 150 141 154 145
rect 145 136 149 140
rect 150 136 154 140
rect 145 131 149 135
rect 150 131 154 135
rect 145 126 149 130
rect 150 126 154 130
rect 145 121 149 125
rect 150 121 154 125
rect 145 116 149 120
rect 150 116 154 120
rect 145 111 149 115
rect 150 111 154 115
rect 203 120 207 124
rect 208 120 212 124
rect 213 120 217 124
rect 218 120 222 124
rect 223 120 227 124
rect 228 120 232 124
rect 233 120 237 124
rect 238 120 242 124
rect 243 120 247 124
rect 248 120 252 124
rect 253 120 257 124
rect 258 120 262 124
rect 263 120 267 124
rect 203 115 207 119
rect 208 115 212 119
rect 213 115 217 119
rect 218 115 222 119
rect 223 115 227 119
rect 228 115 232 119
rect 233 115 237 119
rect 238 115 242 119
rect 243 115 247 119
rect 248 115 252 119
rect 253 115 257 119
rect 258 115 262 119
rect 263 115 267 119
rect 145 106 149 110
rect 150 106 154 110
rect 145 101 149 105
rect 150 101 154 105
rect 145 96 149 100
rect 150 96 154 100
rect 43 63 47 67
rect 48 63 52 67
rect 53 63 57 67
rect 58 63 62 67
rect 63 63 67 67
rect 68 63 72 67
rect 73 63 77 67
rect 78 63 82 67
rect 83 63 87 67
rect 88 63 92 67
rect 93 63 97 67
rect 98 63 102 67
rect 103 63 107 67
rect 43 58 47 62
rect 48 58 52 62
rect 53 58 57 62
rect 58 58 62 62
rect 63 58 67 62
rect 68 58 72 62
rect 73 58 77 62
rect 78 58 82 62
rect 83 58 87 62
rect 88 58 92 62
rect 93 58 97 62
rect 98 58 102 62
rect 103 58 107 62
rect 225 63 229 67
rect 230 63 234 67
rect 235 63 239 67
rect 240 63 244 67
rect 245 63 249 67
rect 250 63 254 67
rect 255 63 259 67
rect 260 63 264 67
rect 265 63 269 67
rect 270 63 274 67
rect 275 63 279 67
rect 225 58 229 62
rect 230 58 234 62
rect 235 58 239 62
rect 240 58 244 62
rect 245 58 249 62
rect 250 58 254 62
rect 255 58 259 62
rect 260 58 264 62
rect 265 58 269 62
rect 270 58 274 62
rect 275 58 279 62
<< metal3 >>
rect 8 155 20 157
rect 8 151 10 155
rect 14 151 15 155
rect 19 151 20 155
rect 8 150 20 151
rect 8 146 10 150
rect 14 146 15 150
rect 19 146 20 150
rect 8 145 20 146
rect 8 141 10 145
rect 14 141 15 145
rect 19 141 20 145
rect 8 140 20 141
rect 8 136 10 140
rect 14 136 15 140
rect 19 136 20 140
rect 8 135 20 136
rect 8 131 10 135
rect 14 131 15 135
rect 19 131 20 135
rect 8 130 20 131
rect 8 126 10 130
rect 14 126 15 130
rect 19 126 20 130
rect 8 125 20 126
rect 8 121 10 125
rect 14 121 15 125
rect 19 121 20 125
rect 8 120 20 121
rect 8 116 10 120
rect 14 116 15 120
rect 19 116 20 120
rect 8 115 20 116
rect 8 111 10 115
rect 14 111 15 115
rect 19 111 20 115
rect 8 110 20 111
rect 8 106 10 110
rect 14 106 15 110
rect 19 106 20 110
rect 8 105 20 106
rect 8 101 10 105
rect 14 101 15 105
rect 19 101 20 105
rect 8 100 20 101
rect 8 96 10 100
rect 14 96 15 100
rect 19 96 20 100
rect 8 95 20 96
rect 8 91 10 95
rect 14 91 15 95
rect 19 91 20 95
rect 144 150 165 151
rect 144 146 145 150
rect 149 146 150 150
rect 154 146 165 150
rect 144 145 165 146
rect 144 141 145 145
rect 149 141 150 145
rect 154 141 165 145
rect 144 140 165 141
rect 144 136 145 140
rect 149 136 150 140
rect 154 136 165 140
rect 144 135 165 136
rect 144 131 145 135
rect 149 131 150 135
rect 154 131 165 135
rect 144 130 165 131
rect 144 126 145 130
rect 149 126 150 130
rect 154 126 165 130
rect 144 125 165 126
rect 144 121 145 125
rect 149 121 150 125
rect 154 121 165 125
rect 144 120 165 121
rect 144 116 145 120
rect 149 116 150 120
rect 154 116 165 120
rect 144 115 165 116
rect 144 111 145 115
rect 149 111 150 115
rect 154 111 165 115
rect 201 124 269 125
rect 201 120 203 124
rect 207 120 208 124
rect 212 120 213 124
rect 217 120 218 124
rect 222 120 223 124
rect 227 120 228 124
rect 232 120 233 124
rect 237 120 238 124
rect 242 120 243 124
rect 247 120 248 124
rect 252 120 253 124
rect 257 120 258 124
rect 262 120 263 124
rect 267 120 269 124
rect 201 119 269 120
rect 201 115 203 119
rect 207 115 208 119
rect 212 115 213 119
rect 217 115 218 119
rect 222 115 223 119
rect 227 115 228 119
rect 232 115 233 119
rect 237 115 238 119
rect 242 115 243 119
rect 247 115 248 119
rect 252 115 253 119
rect 257 115 258 119
rect 262 115 263 119
rect 267 115 269 119
rect 201 112 269 115
rect 144 110 165 111
rect 144 106 145 110
rect 149 106 150 110
rect 154 106 165 110
rect 144 105 165 106
rect 144 101 145 105
rect 149 101 150 105
rect 154 101 165 105
rect 144 100 165 101
rect 144 96 145 100
rect 149 96 150 100
rect 154 96 165 100
rect 144 94 165 96
rect 8 88 20 91
rect 41 67 109 68
rect 41 63 43 67
rect 47 63 48 67
rect 52 63 53 67
rect 57 63 58 67
rect 62 63 63 67
rect 67 63 68 67
rect 72 63 73 67
rect 77 63 78 67
rect 82 63 83 67
rect 87 63 88 67
rect 92 63 93 67
rect 97 63 98 67
rect 102 63 103 67
rect 107 63 109 67
rect 41 62 109 63
rect 41 58 43 62
rect 47 58 48 62
rect 52 58 53 62
rect 57 58 58 62
rect 62 58 63 62
rect 67 58 68 62
rect 72 58 73 62
rect 77 58 78 62
rect 82 58 83 62
rect 87 58 88 62
rect 92 58 93 62
rect 97 58 98 62
rect 102 58 103 62
rect 107 58 109 62
rect 41 55 109 58
rect 224 67 281 69
rect 224 63 225 67
rect 229 63 230 67
rect 234 63 235 67
rect 239 63 240 67
rect 244 63 245 67
rect 249 63 250 67
rect 254 63 255 67
rect 259 63 260 67
rect 264 63 265 67
rect 269 63 270 67
rect 274 63 275 67
rect 279 63 281 67
rect 224 62 281 63
rect 224 58 225 62
rect 229 58 230 62
rect 234 58 235 62
rect 239 58 240 62
rect 244 58 245 62
rect 249 58 250 62
rect 254 58 255 62
rect 259 58 260 62
rect 264 58 265 62
rect 269 58 270 62
rect 274 58 275 62
rect 279 58 281 62
rect 224 56 281 58
use barepad  b
timestamp 1006127261
transform 1 0 9 0 1 -366
box 16 702 276 1014
use ndiode  nd
timestamp 1037203521
transform 1 0 41 0 1 206
box -14 -13 82 128
use pdiode  pd
timestamp 1037203492
transform 1 0 180 0 1 202
box 7 -9 103 132
use barering  br
timestamp 1006127261
transform 1 0 -2 0 1 -12
box 2 -23 311 176
<< labels >>
rlabel metal1 153 210 153 210 1 Vdd!
rlabel metal3 15 94 15 94 1 Vdd!_uq0
rlabel m3contact 17 98 17 98 1 Vdd!0
<< end >>
