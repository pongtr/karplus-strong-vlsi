magic
tech scmos
timestamp 1007670165
<< ntransistor >>
rect 24 7 28 9
rect 39 7 42 15
rect 24 -1 44 1
rect 24 -6 44 -4
<< ptransistor >>
rect -6 12 -3 15
rect 8 7 12 9
rect -18 -1 12 1
rect -18 -6 12 -4
<< ndiffusion >>
rect 39 15 42 16
rect 24 9 28 10
rect 24 6 28 7
rect 39 6 42 7
rect 42 2 44 4
rect 24 1 44 2
rect 24 -4 44 -1
rect 24 -7 44 -6
rect 28 -9 44 -7
<< pdiffusion >>
rect -6 15 -3 16
rect -18 6 -14 8
rect -6 6 -3 12
rect 8 9 12 10
rect 8 6 12 7
rect -18 1 12 2
rect -18 -4 12 -1
rect -18 -7 12 -6
rect -14 -9 12 -7
<< ndcontact >>
rect 38 16 42 20
rect 24 10 28 14
rect 24 2 42 6
rect 24 -11 28 -7
<< pdcontact >>
rect -6 16 -2 20
rect 8 10 12 14
rect -18 2 12 6
rect -18 -11 -14 -7
<< psubstratepcontact >>
rect 47 8 51 21
<< nsubstratencontact >>
rect -18 8 -14 20
<< polysilicon >>
rect 0 15 36 17
rect -8 12 -6 15
rect -3 13 2 15
rect -3 12 -2 13
rect 6 7 8 9
rect 12 7 16 9
rect 34 13 39 15
rect 38 9 39 13
rect 20 7 24 9
rect 28 7 30 9
rect 37 7 39 9
rect 42 7 44 15
rect -20 -1 -18 1
rect 12 -1 24 1
rect 44 -1 46 1
rect -20 -6 -18 -4
rect 12 -6 14 -4
rect 22 -6 24 -4
rect 44 -6 46 -4
<< polycontact >>
rect -2 9 2 13
rect 16 6 20 10
rect 34 9 38 13
<< metal1 >>
rect -2 17 38 20
rect 2 10 8 13
rect 17 10 20 17
rect 28 10 34 13
rect -18 6 -14 8
rect 47 6 51 8
rect 16 -7 19 6
rect 42 3 51 6
rect -14 -10 24 -7
<< labels >>
rlabel pdcontact -17 -10 -17 -10 1 _out
rlabel polysilicon -19 -5 -19 -5 1 _phi0
rlabel polysilicon -19 0 -19 0 1 in
rlabel pdcontact -17 3 -17 3 1 Vdd!
rlabel ndcontact 25 -10 25 -10 1 _out
rlabel polysilicon 23 -5 23 -5 1 phi0
rlabel polysilicon 23 0 23 0 1 in
rlabel pdcontact 3 4 3 4 1 Vdd!
rlabel ndcontact 33 4 33 4 1 GND!
rlabel ndcontact 25 3 25 3 1 GND!
<< end >>
