magic
tech scmos
timestamp 1006127261
<< psubstratepdiff >>
rect 2 87 311 91
rect 2 83 286 87
rect 290 83 291 87
rect 295 83 296 87
rect 300 83 301 87
rect 305 83 311 87
rect 2 77 311 83
rect 2 73 286 77
rect 290 73 291 77
rect 295 73 296 77
rect 300 73 301 77
rect 305 73 311 77
rect 2 67 311 73
rect 2 63 286 67
rect 290 63 291 67
rect 295 63 296 67
rect 300 63 301 67
rect 305 63 311 67
rect 2 57 311 63
rect 2 53 286 57
rect 290 53 291 57
rect 295 53 296 57
rect 300 53 301 57
rect 305 53 311 57
rect 2 51 311 53
<< nsubstratendiff >>
rect 2 133 311 137
rect 2 129 286 133
rect 290 129 291 133
rect 295 129 296 133
rect 300 129 301 133
rect 305 129 311 133
rect 2 123 311 129
rect 2 119 286 123
rect 290 119 291 123
rect 295 119 296 123
rect 300 119 301 123
rect 305 119 311 123
rect 2 113 311 119
rect 2 109 286 113
rect 290 109 291 113
rect 295 109 296 113
rect 300 109 301 113
rect 305 109 311 113
rect 2 103 311 109
rect 2 99 286 103
rect 290 99 291 103
rect 295 99 296 103
rect 300 99 301 103
rect 305 99 311 103
rect 2 97 311 99
<< psubstratepcontact >>
rect 286 83 290 87
rect 291 83 295 87
rect 296 83 300 87
rect 301 83 305 87
rect 286 73 290 77
rect 291 73 295 77
rect 296 73 300 77
rect 301 73 305 77
rect 286 63 290 67
rect 291 63 295 67
rect 296 63 300 67
rect 301 63 305 67
rect 286 53 290 57
rect 291 53 295 57
rect 296 53 300 57
rect 301 53 305 57
<< nsubstratencontact >>
rect 286 129 290 133
rect 291 129 295 133
rect 296 129 300 133
rect 301 129 305 133
rect 286 119 290 123
rect 291 119 295 123
rect 296 119 300 123
rect 301 119 305 123
rect 286 109 290 113
rect 291 109 295 113
rect 296 109 300 113
rect 301 109 305 113
rect 286 99 290 103
rect 291 99 295 103
rect 296 99 300 103
rect 301 99 305 103
<< metal1 >>
rect 290 129 291 133
rect 295 129 296 133
rect 300 129 301 133
rect 286 128 305 129
rect 290 124 291 128
rect 295 124 296 128
rect 300 124 301 128
rect 286 123 305 124
rect 290 119 291 123
rect 295 119 296 123
rect 300 119 301 123
rect 286 118 305 119
rect 290 114 291 118
rect 295 114 296 118
rect 300 114 301 118
rect 286 113 305 114
rect 290 109 291 113
rect 295 109 296 113
rect 300 109 301 113
rect 286 108 305 109
rect 290 104 291 108
rect 295 104 296 108
rect 300 104 301 108
rect 286 103 305 104
rect 290 99 291 103
rect 295 99 296 103
rect 300 99 301 103
rect 290 83 291 87
rect 295 83 296 87
rect 300 83 301 87
rect 286 82 305 83
rect 290 78 291 82
rect 295 78 296 82
rect 300 78 301 82
rect 286 77 305 78
rect 290 73 291 77
rect 295 73 296 77
rect 300 73 301 77
rect 286 72 305 73
rect 290 68 291 72
rect 295 68 296 72
rect 300 68 301 72
rect 286 67 305 68
rect 290 63 291 67
rect 295 63 296 67
rect 300 63 301 67
rect 286 62 305 63
rect 290 58 291 62
rect 295 58 296 62
rect 300 58 301 62
rect 286 57 305 58
rect 290 53 291 57
rect 295 53 296 57
rect 300 53 301 57
<< m2contact >>
rect 286 124 290 128
rect 291 124 295 128
rect 296 124 300 128
rect 301 124 305 128
rect 286 114 290 118
rect 291 114 295 118
rect 296 114 300 118
rect 301 114 305 118
rect 286 104 290 108
rect 291 104 295 108
rect 296 104 300 108
rect 301 104 305 108
rect 286 78 290 82
rect 291 78 295 82
rect 296 78 300 82
rect 301 78 305 82
rect 286 68 290 72
rect 291 68 295 72
rect 296 68 300 72
rect 301 68 305 72
rect 286 58 290 62
rect 291 58 295 62
rect 296 58 300 62
rect 301 58 305 62
<< metal2 >>
rect 290 129 291 133
rect 295 129 296 133
rect 300 129 301 133
rect 286 128 305 129
rect 290 124 291 128
rect 295 124 296 128
rect 300 124 301 128
rect 286 123 305 124
rect 290 119 291 123
rect 295 119 296 123
rect 300 119 301 123
rect 286 118 305 119
rect 290 114 291 118
rect 295 114 296 118
rect 300 114 301 118
rect 286 113 305 114
rect 290 109 291 113
rect 295 109 296 113
rect 300 109 301 113
rect 286 108 305 109
rect 290 104 291 108
rect 295 104 296 108
rect 300 104 301 108
rect 286 103 305 104
rect 290 99 291 103
rect 295 99 296 103
rect 300 99 301 103
rect 290 83 291 87
rect 295 83 296 87
rect 300 83 301 87
rect 286 82 305 83
rect 290 78 291 82
rect 295 78 296 82
rect 300 78 301 82
rect 286 77 305 78
rect 290 73 291 77
rect 295 73 296 77
rect 300 73 301 77
rect 286 72 305 73
rect 290 68 291 72
rect 295 68 296 72
rect 300 68 301 72
rect 286 67 305 68
rect 290 63 291 67
rect 295 63 296 67
rect 300 63 301 67
rect 286 62 305 63
rect 290 58 291 62
rect 295 58 296 62
rect 300 58 301 62
rect 286 57 305 58
rect 290 53 291 57
rect 295 53 296 57
rect 300 53 301 57
<< m3contact >>
rect 286 129 290 133
rect 291 129 295 133
rect 296 129 300 133
rect 301 129 305 133
rect 286 119 290 123
rect 291 119 295 123
rect 296 119 300 123
rect 301 119 305 123
rect 286 109 290 113
rect 291 109 295 113
rect 296 109 300 113
rect 301 109 305 113
rect 286 99 290 103
rect 291 99 295 103
rect 296 99 300 103
rect 301 99 305 103
rect 286 83 290 87
rect 291 83 295 87
rect 296 83 300 87
rect 301 83 305 87
rect 286 73 290 77
rect 291 73 295 77
rect 296 73 300 77
rect 301 73 305 77
rect 286 63 290 67
rect 291 63 295 67
rect 296 63 300 67
rect 301 63 305 67
rect 286 53 290 57
rect 291 53 295 57
rect 296 53 300 57
rect 301 53 305 57
<< metal3 >>
rect 2 133 311 176
rect 2 129 286 133
rect 290 129 291 133
rect 295 129 296 133
rect 300 129 301 133
rect 305 129 311 133
rect 2 123 311 129
rect 2 119 286 123
rect 290 119 291 123
rect 295 119 296 123
rect 300 119 301 123
rect 305 119 311 123
rect 2 113 311 119
rect 2 109 286 113
rect 290 109 291 113
rect 295 109 296 113
rect 300 109 301 113
rect 305 109 311 113
rect 2 103 311 109
rect 2 99 286 103
rect 290 99 291 103
rect 295 99 296 103
rect 300 99 301 103
rect 305 99 311 103
rect 2 96 311 99
rect 2 87 311 92
rect 2 83 286 87
rect 290 83 291 87
rect 295 83 296 87
rect 300 83 301 87
rect 305 83 311 87
rect 2 77 311 83
rect 2 73 286 77
rect 290 73 291 77
rect 295 73 296 77
rect 300 73 301 77
rect 305 73 311 77
rect 2 67 311 73
rect 2 63 286 67
rect 290 63 291 67
rect 295 63 296 67
rect 300 63 301 67
rect 305 63 311 67
rect 2 57 311 63
rect 2 53 286 57
rect 290 53 291 57
rect 295 53 296 57
rect 300 53 301 57
rect 305 53 311 57
rect 2 -23 311 53
<< labels >>
rlabel metal3 16 107 16 107 1 Vdd!
rlabel metal3 15 81 15 81 1 GND!
<< end >>
