magic
tech scmos
timestamp 1006127261
<< nwell >>
rect 16 754 276 1014
<< metal1 >>
rect 16 1011 276 1014
rect 16 757 19 1011
rect 273 757 276 1011
rect 16 754 276 757
rect 58 744 234 754
rect 68 734 224 744
rect 78 724 214 734
rect 88 714 204 724
rect 98 702 194 714
<< metal2 >>
rect 16 1011 276 1014
rect 16 757 19 1011
rect 273 757 276 1011
rect 16 754 276 757
<< pad >>
rect 19 757 273 1011
<< end >>
