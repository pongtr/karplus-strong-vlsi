magic
tech scmos
timestamp 1512379586
<< nwell >>
rect -16 25 164 53
rect -21 -29 0 -5
<< pwell >>
rect -21 -3 167 22
rect 1 -29 166 -3
<< ntransistor >>
rect 1 9 3 16
rect 6 9 8 16
rect 14 9 16 16
rect 19 9 21 16
rect 27 9 29 16
rect 32 9 34 16
rect 44 9 46 16
rect 52 9 54 16
rect 60 9 62 16
rect 68 9 70 16
rect 76 9 78 16
rect 84 9 86 16
rect 92 9 94 16
rect 100 9 102 16
rect 108 9 110 16
rect 116 9 118 16
rect 124 9 126 16
rect 132 9 134 16
rect 9 -6 13 -4
rect 52 -2 54 2
rect 149 6 153 8
rect 21 -18 25 -16
<< ptransistor >>
rect 52 42 54 46
rect 92 43 94 47
rect -5 31 -3 38
rect 3 31 5 38
rect 11 31 13 38
rect 19 31 21 38
rect 27 31 29 38
rect 35 31 37 38
rect 44 31 46 38
rect 51 31 53 38
rect 60 31 62 38
rect 68 31 70 38
rect 76 31 78 38
rect 84 31 86 38
rect 92 31 94 38
rect 100 31 102 38
rect 108 31 110 38
rect 116 31 118 38
rect 124 31 126 38
rect 132 31 134 38
rect 140 31 142 38
rect -10 -18 -6 -16
<< ndiffusion >>
rect 0 9 1 16
rect 3 9 6 16
rect 8 9 14 16
rect 16 9 19 16
rect 21 9 22 16
rect 26 9 27 16
rect 29 9 32 16
rect 34 9 37 16
rect 41 9 44 16
rect 46 13 52 16
rect 46 9 47 13
rect 51 9 52 13
rect 54 12 55 16
rect 59 12 60 16
rect 54 9 60 12
rect 62 13 68 16
rect 62 9 63 13
rect 67 9 68 13
rect 70 12 71 16
rect 75 12 76 16
rect 70 9 76 12
rect 78 13 84 16
rect 78 9 79 13
rect 83 9 84 13
rect 86 12 87 16
rect 91 12 92 16
rect 86 9 92 12
rect 94 13 100 16
rect 94 9 95 13
rect 99 9 100 13
rect 102 12 103 16
rect 107 12 108 16
rect 102 9 108 12
rect 110 13 116 16
rect 110 9 111 13
rect 115 9 116 13
rect 118 12 119 16
rect 123 12 124 16
rect 118 9 124 12
rect 126 13 132 16
rect 126 9 127 13
rect 131 9 132 13
rect 134 9 135 16
rect 9 2 13 9
rect 9 -4 13 -2
rect 9 -9 13 -6
rect 21 -16 25 -2
rect 51 -2 52 2
rect 54 -2 55 2
rect 149 8 153 9
rect 149 5 153 6
rect 21 -19 25 -18
<< pdiffusion >>
rect 42 42 52 46
rect 54 42 55 46
rect 38 38 42 42
rect 91 43 92 47
rect 94 43 95 47
rect -6 31 -5 38
rect -3 31 -2 38
rect 2 31 3 38
rect 5 34 6 38
rect 10 34 11 38
rect 5 31 11 34
rect 13 31 14 38
rect 18 31 19 38
rect 21 31 22 38
rect 26 31 27 38
rect 29 31 30 38
rect 34 31 35 38
rect 37 31 44 38
rect 46 31 51 38
rect 53 31 60 38
rect 62 31 63 38
rect 67 31 68 38
rect 70 31 76 38
rect 78 31 84 38
rect 86 34 87 38
rect 91 34 92 38
rect 86 31 92 34
rect 94 31 100 38
rect 102 31 108 38
rect 110 31 111 38
rect 115 31 116 38
rect 118 31 124 38
rect 126 31 132 38
rect 134 31 135 38
rect 139 31 140 38
rect 142 31 143 38
rect -10 -16 -6 -15
rect -10 -19 -6 -18
<< ndcontact >>
rect -4 9 0 16
rect 22 9 26 16
rect 37 9 41 16
rect 47 9 51 13
rect 55 12 59 16
rect 63 9 67 13
rect 71 12 75 16
rect 79 9 83 13
rect 87 12 91 16
rect 95 9 99 13
rect 103 12 107 16
rect 111 9 115 13
rect 119 12 123 16
rect 127 9 131 13
rect 135 9 139 16
rect 9 -2 13 2
rect 21 -2 25 2
rect 9 -13 13 -9
rect 47 -2 51 2
rect 55 -2 59 2
rect 149 9 153 13
rect 149 1 153 5
rect 21 -23 25 -19
<< pdcontact >>
rect 38 42 42 46
rect 55 42 59 46
rect 87 43 91 47
rect 95 43 99 47
rect -10 31 -6 38
rect -2 31 2 38
rect 6 34 10 38
rect 14 31 18 38
rect 22 31 26 38
rect 30 31 34 38
rect 63 31 67 38
rect 87 34 91 38
rect 111 31 115 38
rect 135 31 139 38
rect 143 31 147 38
rect -10 -15 -6 -11
rect -10 -23 -6 -19
<< nsubstratendiff >>
rect -18 -26 -14 -25
<< psubstratepcontact >>
rect -14 11 -10 15
<< nsubstratencontact >>
rect 156 33 160 37
rect -18 -25 -14 -21
<< polysilicon >>
rect -27 71 102 73
rect -27 62 -3 64
rect -5 55 -3 62
rect -5 53 86 55
rect -5 38 -3 53
rect 11 48 54 50
rect 3 38 5 40
rect 11 38 13 48
rect 19 38 21 40
rect 27 38 29 40
rect 35 38 37 48
rect 52 46 54 48
rect 52 41 54 42
rect 44 38 46 41
rect 51 39 54 41
rect 51 38 53 39
rect 60 38 62 40
rect 68 38 70 40
rect 76 38 78 42
rect 84 38 86 53
rect 92 47 94 49
rect 92 38 94 43
rect 100 38 102 71
rect 108 38 110 40
rect 116 38 118 40
rect 124 38 126 40
rect 132 38 134 47
rect 140 38 142 40
rect -5 28 -3 31
rect 3 28 5 31
rect -5 26 5 28
rect 1 16 3 26
rect 11 21 13 31
rect 19 28 21 31
rect 27 28 29 31
rect 35 29 37 31
rect 19 24 22 28
rect 26 24 29 28
rect 6 19 16 21
rect 6 16 8 19
rect 14 16 16 19
rect 19 16 21 24
rect 27 16 29 24
rect 32 16 34 18
rect 44 16 46 31
rect 51 20 53 31
rect 60 21 62 31
rect 68 21 70 31
rect 51 17 54 20
rect 52 16 54 17
rect 60 19 70 21
rect 60 16 62 19
rect 68 16 70 19
rect 76 16 78 31
rect 84 29 86 31
rect 92 29 94 31
rect 84 27 94 29
rect 84 16 86 27
rect 92 16 94 27
rect 100 16 102 31
rect 108 16 110 31
rect 116 16 118 31
rect 124 16 126 31
rect 132 16 134 31
rect 1 -4 3 9
rect 6 7 8 9
rect 14 7 16 9
rect 19 7 21 9
rect 1 -6 9 -4
rect 13 -5 20 -4
rect 13 -6 16 -5
rect 27 -16 29 9
rect 32 -5 34 9
rect 44 -13 46 9
rect 52 2 54 9
rect 60 7 62 9
rect 68 7 70 9
rect 76 2 78 9
rect 84 7 86 9
rect 92 7 94 9
rect 52 -6 54 -2
rect 100 -6 102 9
rect 108 7 110 9
rect 116 7 118 9
rect 108 5 118 7
rect 116 -6 118 5
rect 124 2 126 9
rect 52 -8 102 -6
rect 132 -13 134 9
rect 140 8 142 31
rect 140 6 149 8
rect 153 6 155 8
rect 143 1 145 6
rect 44 -15 134 -13
rect -12 -18 -10 -16
rect -6 -18 21 -16
rect 25 -18 29 -16
<< polycontact >>
rect 75 42 79 46
rect 128 43 132 47
rect 22 24 26 28
rect 56 24 60 28
rect 16 -9 20 -5
rect 32 -9 36 -5
rect 40 -16 44 -12
rect 75 -2 79 2
rect 123 -2 127 2
rect 115 -10 119 -6
rect 142 -3 146 1
<< metal1 >>
rect -27 53 167 56
rect -10 38 -6 53
rect -2 47 34 50
rect -2 38 2 47
rect 6 41 26 44
rect 6 38 10 41
rect 22 38 26 41
rect 30 38 34 47
rect 38 46 42 53
rect 87 47 91 53
rect 59 42 75 46
rect 99 43 128 47
rect 87 38 91 43
rect 135 38 139 53
rect -25 -35 -21 20
rect -10 -7 -7 31
rect 14 28 18 31
rect 63 30 67 31
rect 111 30 115 31
rect -4 25 18 28
rect -4 16 0 25
rect 26 24 56 28
rect 63 27 123 30
rect 119 20 123 27
rect 143 24 147 31
rect 143 20 163 24
rect 37 17 59 20
rect 37 16 41 17
rect -4 8 0 9
rect 55 16 59 17
rect 22 8 26 9
rect -4 5 26 8
rect 37 2 41 9
rect 71 17 107 20
rect 71 16 75 17
rect 47 8 51 9
rect 87 16 91 17
rect 63 8 67 9
rect 103 16 107 17
rect 79 8 83 9
rect 47 5 83 8
rect 119 17 139 20
rect 119 16 123 17
rect 95 8 99 9
rect 135 16 139 17
rect 111 8 115 9
rect 127 8 131 9
rect 95 5 131 8
rect 143 13 147 20
rect 143 9 149 13
rect 13 -2 21 2
rect 25 -2 47 2
rect 59 -2 75 2
rect 79 -2 123 2
rect -10 -11 -6 -7
rect 20 -9 32 -5
rect 13 -13 40 -12
rect 9 -16 40 -13
rect 115 -19 119 -10
rect -6 -23 21 -19
rect 25 -23 119 -19
rect 135 -17 139 9
rect 149 5 153 6
rect 135 -21 169 -17
rect -10 -32 -6 -23
<< m2contact >>
rect -25 20 -21 24
rect 22 20 26 24
rect 156 29 160 33
rect 163 20 167 24
rect 26 5 30 9
rect 5 -2 9 2
rect -18 -29 -14 -25
rect 149 -3 153 1
rect 142 -7 146 -3
rect -25 -39 -21 -35
<< metal2 >>
rect -21 20 22 24
rect -27 -29 -18 -26
rect 5 -26 9 -2
rect 30 -4 33 9
rect 30 -7 142 -4
rect 149 -26 153 -3
rect 156 -26 160 29
rect 163 24 167 85
rect -14 -29 169 -26
rect -21 -39 169 -35
<< labels >>
rlabel metal2 -13 22 -13 22 3 cin
rlabel polysilicon -4 57 -4 57 5 a
rlabel polysilicon 101 57 101 57 5 b
rlabel metal1 -13 54 -13 54 4 Vdd!
rlabel metal1 63 0 63 0 1 _b
rlabel metal1 16 27 16 27 1 _cout
rlabel metal2 -11 -28 -11 -28 2 GND!
rlabel metal1 31 -21 31 -21 1 _cin
rlabel metal1 13 -14 13 -14 1 _a
rlabel metal1 151 22 151 22 1 cout
rlabel metal1 168 -21 168 -17 7 s
<< end >>
