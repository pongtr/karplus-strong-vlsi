magic
tech scmos
timestamp 1512633651
use latch_one  latch_one_0
array 0 0 142 0 10 124
timestamp 1512631377
transform 1 0 49 0 1 -1217
box -49 1249 93 1373
<< end >>
