magic
tech scmos
timestamp 1512361937
use sreg_10b  sreg_10b_0
array 0 63 56 0 0 1248
timestamp 1512361937
transform 1 0 0 0 1 3
box 0 -3 56 1245
<< end >>
