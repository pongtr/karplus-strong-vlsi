magic
tech scmos
timestamp 1508969492
<< checkpaint >>
rect -1 -270 365 34
<< polysilicon >>
rect 308 21 315 23
rect 319 21 323 23
rect 327 21 331 23
rect 335 21 339 23
rect 343 21 350 23
rect 10 -2 12 3
rect 10 -10 12 -6
rect 10 -18 12 -14
rect 10 -26 12 -22
rect 10 -34 12 -30
rect 34 -34 36 8
rect 42 -2 44 8
rect 42 -10 44 -6
rect 10 -42 12 -38
rect 34 -42 36 -38
rect 10 -51 12 -46
rect 34 -56 36 -46
rect 42 -56 44 -14
rect 50 -26 52 8
rect 58 -2 60 8
rect 58 -10 60 -6
rect 66 -10 68 8
rect 74 -2 76 8
rect 58 -18 60 -14
rect 66 -18 68 -14
rect 50 -42 52 -30
rect 58 -34 60 -22
rect 50 -56 52 -46
rect 58 -56 60 -38
rect 66 -56 68 -22
rect 74 -26 76 -6
rect 82 -18 84 8
rect 74 -34 76 -30
rect 82 -34 84 -22
rect 90 -26 92 8
rect 111 5 113 7
rect 117 5 129 7
rect 133 5 136 7
rect 140 5 169 7
rect 173 5 185 7
rect 189 5 191 7
rect 103 -3 113 -1
rect 117 -3 140 -1
rect 144 -3 146 -1
rect 207 0 238 2
rect 258 0 270 2
rect 280 0 282 2
rect 158 -3 161 -1
rect 165 -3 185 -1
rect 189 -3 191 -1
rect 103 -12 105 -3
rect 111 -11 113 -9
rect 117 -11 129 -9
rect 133 -11 136 -9
rect 310 -3 315 -1
rect 319 -3 355 -1
rect 207 -8 208 -6
rect 228 -8 290 -6
rect 300 -8 302 -6
rect 140 -11 169 -9
rect 173 -11 185 -9
rect 189 -11 191 -9
rect 103 -19 113 -17
rect 117 -19 140 -17
rect 144 -19 146 -17
rect 310 -11 331 -9
rect 335 -11 355 -9
rect 207 -16 238 -14
rect 258 -16 270 -14
rect 280 -16 282 -14
rect 158 -19 161 -17
rect 165 -19 185 -17
rect 189 -19 191 -17
rect 103 -28 105 -19
rect 111 -27 113 -25
rect 117 -27 129 -25
rect 133 -27 136 -25
rect 74 -42 76 -38
rect 74 -56 76 -46
rect 82 -56 84 -38
rect 90 -42 92 -30
rect 310 -19 339 -17
rect 343 -19 355 -17
rect 207 -24 208 -22
rect 228 -24 290 -22
rect 300 -24 302 -22
rect 140 -27 169 -25
rect 173 -27 185 -25
rect 189 -27 191 -25
rect 103 -35 113 -33
rect 117 -35 140 -33
rect 144 -35 146 -33
rect 310 -27 315 -25
rect 319 -27 355 -25
rect 207 -32 238 -30
rect 258 -32 270 -30
rect 280 -32 282 -30
rect 158 -35 161 -33
rect 165 -35 185 -33
rect 189 -35 191 -33
rect 103 -44 105 -35
rect 310 -35 323 -33
rect 327 -35 355 -33
rect 207 -40 208 -38
rect 228 -40 290 -38
rect 300 -40 302 -38
rect 310 -43 323 -41
rect 327 -43 355 -41
rect 90 -56 92 -46
rect 327 -54 330 -52
rect 343 -54 346 -52
rect 328 -64 330 -54
rect 40 -66 42 -64
rect 56 -66 58 -64
rect 72 -66 74 -64
rect 88 -66 90 -64
rect 32 -89 34 -87
rect 32 -114 34 -102
rect 32 -176 34 -139
rect 40 -149 42 -79
rect 48 -89 50 -87
rect 48 -114 50 -102
rect 40 -176 42 -175
rect 48 -176 50 -139
rect 56 -149 58 -79
rect 64 -89 66 -87
rect 64 -114 66 -102
rect 56 -176 58 -175
rect 64 -176 66 -139
rect 72 -149 74 -79
rect 344 -64 346 -54
rect 320 -79 322 -78
rect 80 -89 82 -87
rect 80 -114 82 -102
rect 72 -176 74 -175
rect 80 -176 82 -139
rect 88 -149 90 -79
rect 320 -93 322 -89
rect 320 -101 322 -99
rect 320 -126 322 -125
rect 328 -128 330 -76
rect 336 -79 338 -78
rect 336 -93 338 -89
rect 336 -101 338 -99
rect 336 -126 338 -125
rect 88 -176 90 -175
rect 39 -192 41 -191
rect 36 -193 41 -192
rect 45 -193 47 -191
rect 55 -192 57 -191
rect 52 -193 57 -192
rect 61 -193 63 -191
rect 71 -192 73 -191
rect 68 -193 73 -192
rect 77 -193 79 -191
rect 87 -192 89 -191
rect 84 -193 89 -192
rect 93 -193 95 -191
rect 38 -198 41 -196
rect 45 -198 47 -196
rect 54 -198 57 -196
rect 61 -198 63 -196
rect 70 -198 73 -196
rect 77 -198 79 -196
rect 86 -198 89 -196
rect 93 -198 95 -196
rect 320 -197 322 -130
rect 344 -128 346 -76
rect 328 -154 330 -152
rect 328 -169 330 -166
rect 38 -206 40 -198
rect 54 -206 56 -198
rect 70 -206 72 -198
rect 86 -206 88 -198
rect 39 -224 41 -223
rect 36 -225 41 -224
rect 45 -225 47 -223
rect 55 -224 57 -223
rect 52 -225 57 -224
rect 61 -225 63 -223
rect 71 -224 73 -223
rect 68 -225 73 -224
rect 77 -225 79 -223
rect 320 -223 322 -219
rect 87 -224 89 -223
rect 84 -225 89 -224
rect 93 -225 95 -223
rect 38 -230 41 -228
rect 45 -230 47 -228
rect 54 -230 57 -228
rect 61 -230 63 -228
rect 70 -230 73 -228
rect 77 -230 79 -228
rect 86 -230 89 -228
rect 93 -230 95 -228
rect 38 -240 40 -230
rect 54 -240 56 -230
rect 70 -240 72 -230
rect 86 -240 88 -230
rect 320 -231 322 -229
rect 320 -244 322 -243
rect 38 -252 40 -244
rect 54 -252 56 -244
rect 70 -252 72 -244
rect 86 -252 88 -244
rect 328 -246 330 -193
rect 336 -197 338 -130
rect 344 -154 346 -152
rect 344 -169 346 -166
rect 336 -223 338 -219
rect 336 -231 338 -229
rect 336 -244 338 -243
rect 38 -254 41 -252
rect 45 -254 47 -252
rect 54 -254 57 -252
rect 61 -254 63 -252
rect 70 -254 73 -252
rect 77 -254 79 -252
rect 86 -254 89 -252
rect 93 -254 95 -252
rect 37 -258 41 -257
rect 39 -259 41 -258
rect 45 -259 47 -257
rect 53 -258 57 -257
rect 55 -259 57 -258
rect 61 -259 63 -257
rect 69 -258 73 -257
rect 71 -259 73 -258
rect 77 -259 79 -257
rect 85 -258 89 -257
rect 87 -259 89 -258
rect 93 -259 95 -257
rect 344 -246 346 -193
rect 328 -260 330 -258
rect 344 -260 346 -258
<< ndiffusion >>
rect 37 -2 41 1
rect 37 -6 42 -2
rect 44 -6 45 -2
rect 37 -10 41 -6
rect 37 -14 42 -10
rect 44 -14 45 -10
rect 37 -34 41 -14
rect 33 -38 34 -34
rect 36 -38 41 -34
rect 37 -42 41 -38
rect 33 -46 34 -42
rect 36 -46 41 -42
rect 37 -49 41 -46
rect 53 -2 57 1
rect 53 -6 58 -2
rect 60 -6 61 -2
rect 53 -10 57 -6
rect 69 -2 73 1
rect 69 -6 74 -2
rect 76 -6 77 -2
rect 69 -10 73 -6
rect 53 -14 58 -10
rect 60 -14 61 -10
rect 65 -14 66 -10
rect 68 -14 73 -10
rect 53 -18 57 -14
rect 69 -18 73 -14
rect 53 -22 58 -18
rect 60 -22 61 -18
rect 65 -22 66 -18
rect 68 -22 73 -18
rect 53 -26 57 -22
rect 49 -30 50 -26
rect 52 -30 57 -26
rect 53 -34 57 -30
rect 53 -38 58 -34
rect 60 -38 61 -34
rect 53 -42 57 -38
rect 49 -46 50 -42
rect 52 -46 57 -42
rect 53 -49 57 -46
rect 69 -26 73 -22
rect 85 -18 89 1
rect 81 -22 82 -18
rect 84 -22 89 -18
rect 69 -30 74 -26
rect 76 -30 77 -26
rect 69 -34 73 -30
rect 85 -26 89 -22
rect 129 7 133 8
rect 129 3 133 5
rect 169 7 173 8
rect 169 3 173 5
rect 129 0 144 3
rect 140 -1 144 0
rect 161 0 173 3
rect 161 -1 165 0
rect 270 2 280 3
rect 140 -4 144 -3
rect 161 -4 165 -3
rect 140 -7 143 -4
rect 129 -9 133 -8
rect 129 -13 133 -11
rect 169 -9 173 -8
rect 270 -1 280 0
rect 315 -1 319 0
rect 282 -5 283 -1
rect 287 -5 288 -1
rect 298 -5 300 -1
rect 315 -4 319 -3
rect 290 -6 300 -5
rect 311 -8 348 -4
rect 290 -9 300 -8
rect 331 -9 335 -8
rect 169 -13 173 -11
rect 129 -16 144 -13
rect 140 -17 144 -16
rect 161 -16 173 -13
rect 161 -17 165 -16
rect 331 -12 335 -11
rect 270 -14 280 -13
rect 85 -30 90 -26
rect 92 -30 93 -26
rect 140 -20 144 -19
rect 161 -20 165 -19
rect 140 -23 143 -20
rect 129 -25 133 -24
rect 85 -34 89 -30
rect 69 -38 74 -34
rect 76 -38 77 -34
rect 81 -38 82 -34
rect 84 -38 89 -34
rect 69 -42 73 -38
rect 69 -46 74 -42
rect 76 -46 77 -42
rect 69 -49 73 -46
rect 85 -42 89 -38
rect 129 -29 133 -27
rect 169 -25 173 -24
rect 270 -17 280 -16
rect 339 -17 343 -16
rect 282 -21 283 -17
rect 287 -21 288 -17
rect 298 -21 300 -17
rect 339 -20 343 -19
rect 290 -22 300 -21
rect 311 -24 348 -20
rect 290 -25 300 -24
rect 315 -25 319 -24
rect 169 -29 173 -27
rect 129 -32 144 -29
rect 140 -33 144 -32
rect 161 -32 173 -29
rect 161 -33 165 -32
rect 315 -28 319 -27
rect 270 -30 280 -29
rect 85 -46 90 -42
rect 92 -46 93 -42
rect 140 -36 144 -35
rect 161 -36 165 -35
rect 140 -39 143 -36
rect 270 -33 280 -32
rect 323 -33 327 -32
rect 282 -37 283 -33
rect 287 -37 288 -33
rect 298 -37 300 -33
rect 323 -36 327 -35
rect 290 -38 300 -37
rect 311 -40 348 -36
rect 290 -41 300 -40
rect 323 -41 327 -40
rect 323 -44 327 -43
rect 85 -49 89 -46
rect 331 -62 335 -61
rect 37 -68 40 -66
rect 39 -79 40 -68
rect 42 -79 43 -66
rect 53 -68 56 -66
rect 35 -82 39 -81
rect 35 -87 39 -86
rect 31 -102 32 -89
rect 34 -102 35 -89
rect 55 -79 56 -68
rect 58 -79 59 -66
rect 69 -68 72 -66
rect 51 -82 55 -81
rect 51 -87 55 -86
rect 47 -102 48 -89
rect 50 -102 51 -89
rect 71 -79 72 -68
rect 74 -79 75 -66
rect 85 -68 88 -66
rect 67 -82 71 -81
rect 67 -87 71 -86
rect 63 -102 64 -89
rect 66 -102 67 -89
rect 87 -79 88 -68
rect 90 -79 91 -66
rect 324 -76 328 -64
rect 330 -71 331 -64
rect 347 -62 351 -61
rect 330 -76 334 -71
rect 324 -79 327 -76
rect 83 -82 87 -81
rect 83 -87 87 -86
rect 79 -102 80 -89
rect 82 -102 83 -89
rect 316 -81 320 -79
rect 319 -89 320 -81
rect 322 -89 327 -79
rect 340 -76 344 -64
rect 346 -71 347 -64
rect 346 -76 350 -71
rect 340 -79 343 -76
rect 332 -81 336 -79
rect 335 -89 336 -81
rect 338 -89 343 -79
rect 319 -241 320 -231
rect 316 -243 320 -241
rect 322 -243 327 -231
rect 47 -251 48 -247
rect 41 -252 45 -251
rect 63 -251 64 -247
rect 57 -252 61 -251
rect 79 -251 80 -247
rect 73 -252 77 -251
rect 95 -251 96 -247
rect 324 -246 327 -243
rect 335 -241 336 -231
rect 332 -243 336 -241
rect 338 -243 343 -231
rect 89 -252 93 -251
rect 41 -257 45 -254
rect 57 -257 61 -254
rect 73 -257 77 -254
rect 89 -257 93 -254
rect 41 -260 45 -259
rect 41 -263 42 -260
rect 57 -260 61 -259
rect 57 -263 58 -260
rect 73 -260 77 -259
rect 73 -263 74 -260
rect 324 -258 328 -246
rect 330 -251 334 -246
rect 340 -246 343 -243
rect 330 -258 331 -251
rect 89 -260 93 -259
rect 340 -258 344 -246
rect 346 -251 350 -246
rect 346 -258 347 -251
rect 89 -263 90 -260
rect 331 -261 335 -260
rect 347 -261 351 -260
<< pdiffusion >>
rect 313 28 345 29
rect 315 23 319 24
rect 323 23 327 24
rect 331 23 335 24
rect 339 23 343 24
rect 315 20 319 21
rect 323 20 327 21
rect 331 20 335 21
rect 339 20 343 21
rect 110 8 111 12
rect 4 -48 5 0
rect 9 -6 10 -2
rect 12 -6 13 -2
rect 9 -14 10 -10
rect 12 -14 13 -10
rect 9 -22 10 -18
rect 12 -22 13 -18
rect 9 -30 10 -26
rect 12 -30 13 -26
rect 9 -38 10 -34
rect 12 -38 13 -34
rect 9 -46 10 -42
rect 12 -46 13 -42
rect 113 7 117 8
rect 113 4 117 5
rect 191 8 192 12
rect 185 7 189 8
rect 113 -1 117 0
rect 185 4 189 5
rect 238 3 243 7
rect 185 -1 189 0
rect 238 2 258 3
rect 238 -1 258 0
rect 113 -4 117 -3
rect 185 -4 189 -3
rect 110 -8 111 -4
rect 113 -9 117 -8
rect 113 -12 117 -11
rect 191 -8 192 -4
rect 208 -5 210 -1
rect 230 -5 231 -1
rect 235 -5 236 -1
rect 185 -9 189 -8
rect 208 -6 228 -5
rect 208 -9 228 -8
rect 113 -17 117 -16
rect 185 -12 189 -11
rect 208 -13 210 -9
rect 238 -13 243 -9
rect 185 -17 189 -16
rect 238 -14 258 -13
rect 238 -17 258 -16
rect 113 -20 117 -19
rect 185 -20 189 -19
rect 110 -24 111 -20
rect 113 -25 117 -24
rect 113 -28 117 -27
rect 191 -24 192 -20
rect 208 -21 210 -17
rect 230 -21 231 -17
rect 235 -21 236 -17
rect 185 -25 189 -24
rect 208 -22 228 -21
rect 208 -25 228 -24
rect 113 -33 117 -32
rect 185 -28 189 -27
rect 208 -29 210 -25
rect 238 -29 243 -25
rect 185 -33 189 -32
rect 238 -30 258 -29
rect 238 -33 258 -32
rect 113 -36 117 -35
rect 110 -40 111 -36
rect 185 -36 189 -35
rect 191 -40 192 -36
rect 208 -37 210 -33
rect 230 -37 231 -33
rect 235 -37 236 -33
rect 208 -38 228 -37
rect 208 -41 228 -40
rect 208 -45 210 -41
rect 31 -132 32 -114
rect 29 -139 32 -132
rect 34 -139 35 -114
rect 35 -142 39 -141
rect 35 -147 39 -146
rect 47 -132 48 -114
rect 45 -139 48 -132
rect 50 -139 51 -114
rect 39 -173 40 -149
rect 35 -175 40 -173
rect 42 -166 43 -149
rect 42 -175 45 -166
rect 51 -142 55 -141
rect 51 -147 55 -146
rect 63 -132 64 -114
rect 61 -139 64 -132
rect 66 -139 67 -114
rect 55 -173 56 -149
rect 51 -175 56 -173
rect 58 -166 59 -149
rect 58 -175 61 -166
rect 67 -142 71 -141
rect 67 -147 71 -146
rect 79 -132 80 -114
rect 77 -139 80 -132
rect 82 -139 83 -114
rect 71 -173 72 -149
rect 67 -175 72 -173
rect 74 -166 75 -149
rect 74 -175 77 -166
rect 83 -142 87 -141
rect 83 -147 87 -146
rect 319 -123 320 -101
rect 316 -125 320 -123
rect 322 -125 327 -101
rect 324 -128 327 -125
rect 335 -123 336 -101
rect 332 -125 336 -123
rect 338 -125 343 -101
rect 87 -173 88 -149
rect 83 -175 88 -173
rect 90 -166 91 -149
rect 90 -175 93 -166
rect 41 -190 42 -188
rect 41 -191 45 -190
rect 57 -190 58 -188
rect 57 -191 61 -190
rect 73 -190 74 -188
rect 73 -191 77 -190
rect 89 -190 90 -188
rect 89 -191 93 -190
rect 41 -196 45 -193
rect 57 -196 61 -193
rect 73 -196 77 -193
rect 89 -196 93 -193
rect 324 -152 328 -128
rect 330 -133 334 -128
rect 340 -128 343 -125
rect 330 -152 331 -133
rect 331 -155 335 -154
rect 324 -193 328 -169
rect 330 -193 331 -169
rect 324 -197 327 -193
rect 41 -199 45 -198
rect 47 -203 48 -199
rect 57 -199 61 -198
rect 63 -203 64 -199
rect 73 -199 77 -198
rect 79 -203 80 -199
rect 89 -199 93 -198
rect 95 -203 96 -199
rect 41 -222 42 -220
rect 41 -223 45 -222
rect 57 -222 58 -220
rect 57 -223 61 -222
rect 73 -222 74 -220
rect 73 -223 77 -222
rect 89 -222 90 -220
rect 319 -219 320 -197
rect 322 -219 327 -197
rect 89 -223 93 -222
rect 41 -228 45 -225
rect 57 -228 61 -225
rect 73 -228 77 -225
rect 89 -228 93 -225
rect 41 -231 45 -230
rect 47 -235 48 -231
rect 57 -231 61 -230
rect 63 -235 64 -231
rect 73 -231 77 -230
rect 79 -235 80 -231
rect 89 -231 93 -230
rect 95 -235 96 -231
rect 340 -152 344 -128
rect 346 -133 350 -128
rect 346 -152 347 -133
rect 347 -155 351 -154
rect 340 -193 344 -169
rect 346 -193 347 -169
rect 340 -197 343 -193
rect 335 -219 336 -197
rect 338 -219 343 -197
<< metal1 >>
rect 16 26 29 30
rect 97 26 287 32
rect 313 28 345 29
rect 16 24 97 26
rect 16 16 20 24
rect 110 8 111 12
rect 121 8 129 11
rect 137 8 140 12
rect 8 7 12 8
rect 30 2 37 5
rect 41 2 53 5
rect 57 2 69 5
rect 73 2 85 5
rect 89 2 93 5
rect 4 -48 5 0
rect 17 -6 45 -3
rect 49 -6 61 -3
rect 65 -6 77 -3
rect 97 -3 98 -2
rect 81 -6 98 -3
rect 106 -4 110 8
rect 121 4 124 8
rect 117 1 120 4
rect 110 -8 111 -4
rect 121 -8 129 -5
rect 137 -8 140 4
rect 17 -14 45 -11
rect 49 -14 61 -11
rect 97 -11 99 -10
rect 65 -13 99 -11
rect 65 -14 100 -13
rect 17 -22 61 -19
rect 65 -22 77 -19
rect 97 -19 98 -18
rect 81 -22 98 -19
rect 106 -20 110 -8
rect 121 -12 124 -8
rect 117 -15 120 -12
rect 110 -24 111 -20
rect 121 -24 129 -21
rect 137 -24 140 -12
rect 17 -30 45 -27
rect 49 -30 77 -27
rect 81 -30 93 -27
rect 97 -29 99 -26
rect 97 -30 100 -29
rect 17 -38 29 -35
rect 33 -38 61 -35
rect 65 -38 77 -35
rect 97 -35 98 -34
rect 81 -38 98 -35
rect 106 -36 110 -24
rect 121 -28 124 -24
rect 117 -31 120 -28
rect 110 -40 111 -36
rect 17 -46 29 -43
rect 33 -46 45 -43
rect 49 -46 77 -43
rect 81 -46 93 -43
rect 97 -45 99 -42
rect 97 -46 100 -45
rect 106 -48 110 -40
rect 1 -169 5 -48
rect 30 -53 37 -50
rect 41 -53 53 -50
rect 57 -53 69 -50
rect 73 -53 85 -50
rect 89 -53 103 -50
rect 106 -52 115 -48
rect 8 -56 12 -55
rect 100 -60 103 -53
rect 1 -199 5 -173
rect 9 -191 12 -60
rect 35 -61 39 -60
rect 43 -61 47 -60
rect 51 -61 55 -60
rect 59 -61 63 -60
rect 67 -61 71 -60
rect 75 -61 79 -60
rect 83 -61 87 -60
rect 91 -61 95 -60
rect 43 -66 47 -65
rect 59 -66 63 -65
rect 35 -82 39 -81
rect 75 -66 79 -65
rect 51 -82 55 -81
rect 91 -66 95 -65
rect 67 -82 71 -81
rect 107 -68 115 -52
rect 137 -52 140 -28
rect 147 -60 151 26
rect 154 -4 158 -3
rect 161 -4 165 26
rect 192 15 276 19
rect 192 12 196 15
rect 173 8 179 11
rect 191 8 192 12
rect 176 4 179 8
rect 180 1 185 4
rect 192 -4 196 8
rect 236 -1 240 15
rect 283 10 287 26
rect 310 24 313 28
rect 345 24 347 28
rect 302 17 306 20
rect 350 20 354 21
rect 258 4 270 7
rect 261 -1 264 4
rect 283 6 306 10
rect 283 -1 287 6
rect 315 4 318 16
rect 173 -8 179 -5
rect 191 -8 192 -4
rect 230 -5 231 -1
rect 235 -5 236 -1
rect 282 -5 283 -1
rect 287 -5 288 -1
rect 305 -5 306 -1
rect 154 -20 158 -19
rect 161 -20 165 -8
rect 176 -12 179 -8
rect 180 -15 185 -12
rect 192 -20 196 -8
rect 228 -13 229 -9
rect 236 -17 240 -5
rect 258 -12 270 -9
rect 261 -17 264 -12
rect 283 -17 287 -5
rect 300 -13 301 -9
rect 305 -13 306 -9
rect 173 -24 179 -21
rect 191 -24 192 -20
rect 230 -21 231 -17
rect 235 -21 236 -17
rect 282 -21 283 -17
rect 287 -21 288 -17
rect 305 -21 306 -17
rect 154 -36 158 -35
rect 161 -36 165 -24
rect 176 -28 179 -24
rect 180 -31 185 -28
rect 192 -36 196 -24
rect 228 -29 229 -25
rect 236 -33 240 -21
rect 258 -28 270 -25
rect 261 -33 264 -28
rect 283 -33 287 -21
rect 300 -29 301 -25
rect 305 -29 306 -25
rect 315 -28 318 0
rect 323 -28 326 16
rect 331 -12 334 16
rect 339 -12 342 16
rect 348 4 352 6
rect 348 -4 352 0
rect 359 -5 360 -1
rect 348 -12 352 -8
rect 359 -13 360 -9
rect 191 -40 192 -36
rect 230 -37 231 -33
rect 235 -37 236 -33
rect 282 -37 283 -33
rect 287 -37 288 -33
rect 305 -37 306 -33
rect 107 -72 111 -68
rect 83 -82 87 -81
rect 9 -223 12 -195
rect 20 -86 35 -82
rect 39 -86 51 -82
rect 55 -86 67 -82
rect 71 -86 83 -82
rect 87 -86 100 -82
rect 16 -247 20 -86
rect 35 -87 39 -86
rect 51 -87 55 -86
rect 67 -87 71 -86
rect 83 -87 87 -86
rect 27 -107 30 -102
rect 27 -110 35 -107
rect 43 -107 46 -102
rect 43 -110 51 -107
rect 59 -107 62 -102
rect 59 -110 67 -107
rect 75 -107 78 -102
rect 75 -110 83 -107
rect 27 -114 30 -110
rect 43 -114 46 -110
rect 59 -114 62 -110
rect 75 -114 78 -110
rect 91 -114 94 -102
rect 29 -139 35 -135
rect 39 -139 51 -135
rect 35 -142 39 -141
rect 55 -139 67 -135
rect 51 -142 55 -141
rect 71 -139 83 -135
rect 67 -142 71 -141
rect 107 -135 115 -72
rect 87 -139 115 -135
rect 83 -142 87 -141
rect 35 -147 39 -146
rect 29 -173 35 -169
rect 43 -147 47 -146
rect 51 -147 55 -146
rect 39 -173 51 -169
rect 59 -147 63 -146
rect 67 -147 71 -146
rect 55 -173 67 -169
rect 75 -147 79 -146
rect 83 -147 87 -146
rect 71 -173 83 -169
rect 91 -147 95 -146
rect 107 -169 115 -139
rect 87 -173 111 -169
rect 33 -181 37 -180
rect 41 -181 45 -180
rect 49 -181 53 -180
rect 57 -181 61 -180
rect 65 -181 69 -180
rect 73 -181 77 -180
rect 81 -181 85 -180
rect 89 -181 93 -180
rect 42 -186 45 -185
rect 58 -186 61 -185
rect 74 -186 77 -185
rect 90 -186 93 -185
rect 35 -193 39 -192
rect 51 -193 55 -192
rect 67 -193 71 -192
rect 83 -193 87 -192
rect 29 -195 100 -193
rect 26 -196 100 -195
rect 107 -199 115 -173
rect 29 -203 32 -199
rect 36 -203 41 -199
rect 47 -203 48 -199
rect 52 -203 57 -199
rect 63 -203 64 -199
rect 68 -203 73 -199
rect 79 -203 80 -199
rect 84 -203 89 -199
rect 95 -203 96 -199
rect 100 -203 115 -199
rect 41 -210 42 -206
rect 57 -210 58 -206
rect 73 -210 74 -206
rect 89 -210 90 -206
rect 38 -217 45 -214
rect 54 -217 61 -214
rect 70 -217 77 -214
rect 86 -217 93 -214
rect 42 -218 45 -217
rect 58 -218 61 -217
rect 74 -218 77 -217
rect 90 -218 93 -217
rect 35 -225 39 -224
rect 51 -225 55 -224
rect 67 -225 71 -224
rect 83 -225 87 -224
rect 29 -227 100 -225
rect 26 -228 100 -227
rect 107 -231 115 -203
rect 29 -235 32 -231
rect 36 -235 41 -231
rect 47 -235 48 -231
rect 52 -235 57 -231
rect 63 -235 64 -231
rect 68 -235 73 -231
rect 79 -235 80 -231
rect 84 -235 89 -231
rect 95 -235 96 -231
rect 100 -235 115 -231
rect 41 -244 42 -240
rect 57 -244 58 -240
rect 73 -244 74 -240
rect 89 -244 90 -240
rect 16 -251 32 -247
rect 36 -251 41 -247
rect 47 -251 48 -247
rect 52 -251 57 -247
rect 63 -251 64 -247
rect 68 -251 73 -247
rect 79 -251 80 -247
rect 84 -251 89 -247
rect 95 -251 96 -247
rect 29 -257 100 -254
rect 35 -258 39 -257
rect 51 -258 55 -257
rect 67 -258 71 -257
rect 83 -258 87 -257
rect 42 -265 45 -264
rect 58 -265 61 -264
rect 74 -265 77 -264
rect 90 -265 93 -264
rect 38 -268 45 -265
rect 54 -268 61 -265
rect 70 -268 77 -265
rect 86 -268 93 -265
rect 107 -268 115 -235
rect 161 -60 165 -40
rect 119 -254 122 -64
rect 147 -82 151 -64
rect 192 -68 196 -40
rect 228 -45 229 -41
rect 236 -68 240 -37
rect 283 -48 287 -37
rect 300 -45 301 -41
rect 305 -45 306 -41
rect 315 -48 318 -32
rect 323 -44 326 -32
rect 283 -52 291 -48
rect 315 -50 319 -48
rect 323 -50 327 -48
rect 331 -48 334 -16
rect 339 -48 342 -16
rect 348 -20 352 -16
rect 359 -21 360 -17
rect 348 -28 352 -24
rect 359 -29 360 -25
rect 348 -36 352 -32
rect 359 -37 360 -33
rect 348 -44 352 -40
rect 359 -45 360 -41
rect 331 -50 335 -48
rect 339 -50 343 -48
rect 276 -74 279 -56
rect 283 -57 291 -56
rect 283 -60 315 -57
rect 287 -61 315 -60
rect 319 -61 331 -57
rect 335 -61 347 -57
rect 287 -64 291 -61
rect 127 -224 130 -196
rect 119 -268 122 -258
rect 127 -268 130 -228
rect 268 -265 271 -130
rect 276 -245 279 -78
rect 276 -265 279 -249
rect 283 -261 291 -64
rect 331 -62 335 -61
rect 347 -62 351 -61
rect 311 -78 319 -75
rect 323 -78 335 -75
rect 339 -78 351 -75
rect 315 -94 318 -89
rect 331 -94 334 -89
rect 315 -101 318 -98
rect 331 -101 334 -98
rect 311 -130 319 -127
rect 323 -130 335 -127
rect 339 -130 351 -127
rect 331 -155 335 -154
rect 347 -155 351 -154
rect 307 -159 315 -155
rect 319 -159 331 -155
rect 335 -159 347 -155
rect 307 -169 311 -159
rect 327 -166 328 -162
rect 343 -166 344 -162
rect 311 -173 331 -169
rect 335 -173 347 -169
rect 315 -224 318 -219
rect 331 -224 334 -219
rect 315 -231 318 -228
rect 331 -231 334 -228
rect 311 -248 319 -245
rect 323 -248 335 -245
rect 339 -248 351 -245
rect 331 -261 335 -260
rect 347 -261 351 -260
rect 283 -265 315 -261
rect 319 -265 331 -261
rect 335 -265 347 -261
<< metal2 >>
rect 97 23 264 25
rect 9 22 264 23
rect 9 20 101 22
rect 9 12 12 20
rect 9 -56 12 8
rect 16 -82 20 12
rect 26 -49 29 1
rect 34 -54 37 12
rect 42 -54 45 12
rect 50 -54 53 12
rect 58 -54 61 12
rect 66 -54 69 12
rect 74 -54 77 12
rect 82 -54 85 12
rect 90 -54 93 12
rect 261 9 264 22
rect 276 24 306 28
rect 276 19 280 24
rect 302 17 350 20
rect 298 9 301 16
rect 261 6 301 9
rect 310 6 348 10
rect 124 0 165 3
rect 180 0 199 3
rect 102 -4 116 -3
rect 102 -6 154 -4
rect 113 -7 154 -6
rect 162 -5 165 0
rect 265 -4 301 -1
rect 305 -4 360 -1
rect 162 -8 199 -5
rect 124 -16 165 -13
rect 233 -13 301 -10
rect 305 -12 360 -9
rect 180 -16 199 -13
rect 102 -20 116 -19
rect 102 -22 154 -20
rect 113 -23 154 -22
rect 162 -21 165 -16
rect 265 -20 301 -17
rect 305 -20 360 -17
rect 162 -24 199 -21
rect 124 -32 165 -29
rect 233 -29 301 -26
rect 305 -28 360 -25
rect 180 -32 199 -29
rect 102 -36 116 -35
rect 102 -38 154 -36
rect 113 -39 154 -38
rect 162 -37 165 -32
rect 265 -36 301 -33
rect 305 -36 360 -33
rect 162 -40 199 -37
rect 233 -45 301 -42
rect 305 -44 360 -41
rect 34 -57 38 -54
rect 42 -57 46 -54
rect 50 -57 54 -54
rect 58 -57 62 -54
rect 66 -57 70 -54
rect 74 -57 78 -54
rect 82 -57 86 -54
rect 90 -57 94 -54
rect 141 -56 276 -53
rect 35 -61 38 -57
rect 43 -61 46 -57
rect 51 -61 54 -57
rect 59 -61 62 -57
rect 67 -61 70 -57
rect 75 -61 78 -57
rect 83 -61 86 -57
rect 91 -61 94 -57
rect 104 -64 119 -61
rect 151 -64 161 -60
rect 165 -64 283 -60
rect 35 -106 38 -65
rect 43 -142 46 -65
rect 51 -106 54 -65
rect 59 -142 62 -65
rect 67 -106 70 -65
rect 75 -142 78 -65
rect 83 -106 86 -65
rect 91 -142 94 -65
rect 115 -72 192 -68
rect 196 -72 236 -68
rect 280 -78 307 -75
rect 104 -86 147 -82
rect 315 -87 318 -54
rect 331 -87 334 -54
rect 315 -90 327 -87
rect 331 -90 343 -87
rect 272 -130 307 -127
rect 43 -164 46 -146
rect 59 -164 62 -146
rect 75 -164 78 -146
rect 91 -164 94 -146
rect 34 -167 46 -164
rect 50 -167 62 -164
rect 66 -167 78 -164
rect 82 -167 94 -164
rect 5 -173 25 -169
rect 34 -181 37 -167
rect 50 -181 53 -167
rect 66 -181 69 -167
rect 82 -181 85 -167
rect 115 -173 307 -169
rect 41 -189 44 -185
rect 57 -189 60 -185
rect 73 -189 76 -185
rect 89 -189 92 -185
rect 12 -195 25 -192
rect 34 -192 44 -189
rect 50 -192 60 -189
rect 66 -192 76 -189
rect 82 -192 92 -189
rect 5 -203 25 -199
rect 34 -213 37 -192
rect 12 -227 25 -224
rect 34 -265 37 -217
rect 42 -240 45 -210
rect 50 -213 53 -192
rect 42 -268 45 -244
rect 50 -265 53 -217
rect 58 -240 61 -210
rect 66 -213 69 -192
rect 58 -268 61 -244
rect 66 -265 69 -217
rect 74 -240 77 -210
rect 82 -213 85 -192
rect 104 -196 126 -193
rect 315 -197 318 -98
rect 324 -162 327 -90
rect 331 -197 334 -98
rect 340 -162 343 -90
rect 315 -200 326 -197
rect 331 -200 342 -197
rect 74 -268 77 -244
rect 82 -265 85 -217
rect 90 -240 93 -210
rect 104 -228 126 -225
rect 90 -268 93 -244
rect 280 -248 307 -245
rect 104 -257 119 -254
rect 315 -265 318 -228
rect 323 -265 326 -200
rect 331 -265 334 -228
rect 339 -265 342 -200
<< ntransistor >>
rect 42 -6 44 -2
rect 42 -14 44 -10
rect 34 -38 36 -34
rect 34 -46 36 -42
rect 58 -6 60 -2
rect 74 -6 76 -2
rect 58 -14 60 -10
rect 66 -14 68 -10
rect 58 -22 60 -18
rect 66 -22 68 -18
rect 50 -30 52 -26
rect 58 -38 60 -34
rect 50 -46 52 -42
rect 82 -22 84 -18
rect 74 -30 76 -26
rect 129 5 133 7
rect 169 5 173 7
rect 140 -3 144 -1
rect 270 0 280 2
rect 161 -3 165 -1
rect 129 -11 133 -9
rect 315 -3 319 -1
rect 290 -8 300 -6
rect 169 -11 173 -9
rect 140 -19 144 -17
rect 331 -11 335 -9
rect 270 -16 280 -14
rect 161 -19 165 -17
rect 90 -30 92 -26
rect 129 -27 133 -25
rect 74 -38 76 -34
rect 82 -38 84 -34
rect 74 -46 76 -42
rect 339 -19 343 -17
rect 290 -24 300 -22
rect 169 -27 173 -25
rect 140 -35 144 -33
rect 315 -27 319 -25
rect 270 -32 280 -30
rect 161 -35 165 -33
rect 90 -46 92 -42
rect 323 -35 327 -33
rect 290 -40 300 -38
rect 323 -43 327 -41
rect 40 -79 42 -66
rect 32 -102 34 -89
rect 56 -79 58 -66
rect 48 -102 50 -89
rect 72 -79 74 -66
rect 64 -102 66 -89
rect 88 -79 90 -66
rect 328 -76 330 -64
rect 80 -102 82 -89
rect 320 -89 322 -79
rect 344 -76 346 -64
rect 336 -89 338 -79
rect 320 -243 322 -231
rect 336 -243 338 -231
rect 41 -254 45 -252
rect 57 -254 61 -252
rect 73 -254 77 -252
rect 89 -254 93 -252
rect 41 -259 45 -257
rect 57 -259 61 -257
rect 73 -259 77 -257
rect 89 -259 93 -257
rect 328 -258 330 -246
rect 344 -258 346 -246
<< ptransistor >>
rect 315 21 319 23
rect 323 21 327 23
rect 331 21 335 23
rect 339 21 343 23
rect 10 -6 12 -2
rect 10 -14 12 -10
rect 10 -22 12 -18
rect 10 -30 12 -26
rect 10 -38 12 -34
rect 10 -46 12 -42
rect 113 5 117 7
rect 185 5 189 7
rect 113 -3 117 -1
rect 238 0 258 2
rect 185 -3 189 -1
rect 113 -11 117 -9
rect 208 -8 228 -6
rect 185 -11 189 -9
rect 113 -19 117 -17
rect 238 -16 258 -14
rect 185 -19 189 -17
rect 113 -27 117 -25
rect 208 -24 228 -22
rect 185 -27 189 -25
rect 113 -35 117 -33
rect 238 -32 258 -30
rect 185 -35 189 -33
rect 208 -40 228 -38
rect 32 -139 34 -114
rect 48 -139 50 -114
rect 40 -175 42 -149
rect 64 -139 66 -114
rect 56 -175 58 -149
rect 80 -139 82 -114
rect 72 -175 74 -149
rect 320 -125 322 -101
rect 336 -125 338 -101
rect 88 -175 90 -149
rect 41 -193 45 -191
rect 57 -193 61 -191
rect 73 -193 77 -191
rect 89 -193 93 -191
rect 41 -198 45 -196
rect 57 -198 61 -196
rect 73 -198 77 -196
rect 89 -198 93 -196
rect 328 -152 330 -128
rect 328 -193 330 -169
rect 41 -225 45 -223
rect 57 -225 61 -223
rect 73 -225 77 -223
rect 320 -219 322 -197
rect 89 -225 93 -223
rect 41 -230 45 -228
rect 57 -230 61 -228
rect 73 -230 77 -228
rect 89 -230 93 -228
rect 344 -152 346 -128
rect 344 -193 346 -169
rect 336 -219 338 -197
<< polycontact >>
rect 350 21 354 25
rect 306 17 310 21
rect 34 8 38 12
rect 42 8 46 12
rect 50 8 54 12
rect 58 8 62 12
rect 66 8 70 12
rect 74 8 78 12
rect 82 8 86 12
rect 90 8 94 12
rect 8 3 12 7
rect 8 -55 12 -51
rect 136 4 140 8
rect 154 -3 158 1
rect 203 -1 207 3
rect 99 -13 103 -9
rect 136 -12 140 -8
rect 306 -5 310 -1
rect 203 -9 207 -5
rect 355 -5 359 -1
rect 154 -19 158 -15
rect 203 -17 207 -13
rect 306 -13 310 -9
rect 355 -13 359 -9
rect 99 -29 103 -25
rect 136 -28 140 -24
rect 306 -21 310 -17
rect 203 -25 207 -21
rect 355 -21 359 -17
rect 154 -35 158 -31
rect 203 -33 207 -29
rect 306 -29 310 -25
rect 355 -29 359 -25
rect 99 -45 103 -41
rect 306 -37 310 -33
rect 203 -41 207 -37
rect 355 -37 359 -33
rect 306 -45 310 -41
rect 355 -45 359 -41
rect 323 -54 327 -50
rect 339 -54 343 -50
rect 34 -60 38 -56
rect 42 -60 46 -56
rect 50 -60 54 -56
rect 58 -60 62 -56
rect 66 -60 70 -56
rect 74 -60 78 -56
rect 82 -60 86 -56
rect 90 -60 94 -56
rect 319 -78 323 -74
rect 319 -130 323 -126
rect 335 -78 339 -74
rect 32 -180 36 -176
rect 40 -180 44 -176
rect 48 -180 52 -176
rect 56 -180 60 -176
rect 64 -180 68 -176
rect 72 -180 76 -176
rect 80 -180 84 -176
rect 88 -180 92 -176
rect 35 -192 39 -188
rect 51 -192 55 -188
rect 67 -192 71 -188
rect 83 -192 87 -188
rect 335 -130 339 -126
rect 328 -166 332 -162
rect 37 -210 41 -206
rect 53 -210 57 -206
rect 69 -210 73 -206
rect 85 -210 89 -206
rect 35 -224 39 -220
rect 51 -224 55 -220
rect 67 -224 71 -220
rect 83 -224 87 -220
rect 37 -244 41 -240
rect 53 -244 57 -240
rect 69 -244 73 -240
rect 85 -244 89 -240
rect 319 -248 323 -244
rect 344 -166 348 -162
rect 35 -262 39 -258
rect 51 -262 55 -258
rect 67 -262 71 -258
rect 83 -262 87 -258
rect 335 -248 339 -244
<< ndcontact >>
rect 37 1 41 5
rect 45 -6 49 -2
rect 45 -14 49 -10
rect 29 -38 33 -34
rect 29 -46 33 -42
rect 37 -53 41 -49
rect 53 1 57 5
rect 61 -6 65 -2
rect 69 1 73 5
rect 77 -6 81 -2
rect 61 -14 65 -10
rect 61 -22 65 -18
rect 45 -30 49 -26
rect 61 -38 65 -34
rect 45 -46 49 -42
rect 53 -53 57 -49
rect 85 1 89 5
rect 77 -22 81 -18
rect 77 -30 81 -26
rect 129 8 133 12
rect 169 8 173 12
rect 270 3 280 7
rect 315 0 319 4
rect 129 -8 133 -4
rect 143 -8 147 -4
rect 161 -8 165 -4
rect 169 -8 173 -4
rect 270 -5 282 -1
rect 288 -5 298 -1
rect 348 -8 352 -4
rect 270 -13 280 -9
rect 290 -13 300 -9
rect 331 -16 335 -12
rect 339 -16 343 -12
rect 93 -30 97 -26
rect 129 -24 133 -20
rect 143 -24 147 -20
rect 161 -24 165 -20
rect 169 -24 173 -20
rect 77 -38 81 -34
rect 77 -46 81 -42
rect 69 -53 73 -49
rect 270 -21 282 -17
rect 288 -21 298 -17
rect 348 -24 352 -20
rect 270 -29 280 -25
rect 290 -29 300 -25
rect 315 -32 319 -28
rect 323 -32 327 -28
rect 93 -46 97 -42
rect 143 -40 147 -36
rect 161 -40 165 -36
rect 270 -37 282 -33
rect 288 -37 298 -33
rect 348 -40 352 -36
rect 290 -45 300 -41
rect 85 -53 89 -49
rect 323 -48 327 -44
rect 35 -81 39 -68
rect 43 -79 47 -66
rect 27 -102 31 -89
rect 35 -102 39 -87
rect 51 -81 55 -68
rect 59 -79 63 -66
rect 43 -102 47 -89
rect 51 -102 55 -87
rect 67 -81 71 -68
rect 75 -79 79 -66
rect 59 -102 63 -89
rect 67 -102 71 -87
rect 83 -81 87 -68
rect 91 -79 95 -66
rect 331 -71 335 -62
rect 75 -102 79 -89
rect 83 -102 87 -87
rect 315 -89 319 -81
rect 91 -102 95 -89
rect 347 -71 351 -62
rect 331 -89 335 -81
rect 315 -241 319 -231
rect 41 -251 47 -247
rect 57 -251 63 -247
rect 73 -251 79 -247
rect 89 -251 95 -247
rect 331 -241 335 -231
rect 42 -264 46 -260
rect 58 -264 62 -260
rect 74 -264 78 -260
rect 331 -260 335 -251
rect 347 -260 351 -251
rect 90 -264 94 -260
<< pdcontact >>
rect 313 24 345 28
rect 315 16 319 20
rect 323 16 327 20
rect 331 16 335 20
rect 339 16 343 20
rect 111 8 117 12
rect 5 -48 9 0
rect 13 -6 17 -2
rect 13 -14 17 -10
rect 13 -22 17 -18
rect 13 -30 17 -26
rect 13 -38 17 -34
rect 13 -46 17 -42
rect 113 0 117 4
rect 185 8 191 12
rect 185 0 189 4
rect 243 3 258 7
rect 111 -8 117 -4
rect 113 -16 117 -12
rect 185 -8 191 -4
rect 210 -5 230 -1
rect 236 -5 258 -1
rect 185 -16 189 -12
rect 210 -13 228 -9
rect 243 -13 258 -9
rect 111 -24 117 -20
rect 113 -32 117 -28
rect 185 -24 191 -20
rect 210 -21 230 -17
rect 236 -21 258 -17
rect 185 -32 189 -28
rect 210 -29 228 -25
rect 243 -29 258 -25
rect 111 -40 117 -36
rect 185 -40 191 -36
rect 210 -37 230 -33
rect 236 -37 258 -33
rect 210 -45 228 -41
rect 27 -132 31 -114
rect 35 -141 39 -114
rect 35 -173 39 -147
rect 43 -132 47 -114
rect 43 -166 47 -147
rect 51 -141 55 -114
rect 51 -173 55 -147
rect 59 -132 63 -114
rect 59 -166 63 -147
rect 67 -141 71 -114
rect 67 -173 71 -147
rect 75 -132 79 -114
rect 75 -166 79 -147
rect 83 -141 87 -114
rect 83 -173 87 -147
rect 91 -132 95 -114
rect 315 -123 319 -101
rect 331 -123 335 -101
rect 91 -166 95 -147
rect 42 -190 46 -186
rect 58 -190 62 -186
rect 74 -190 78 -186
rect 90 -190 94 -186
rect 331 -154 335 -133
rect 331 -193 335 -169
rect 41 -203 47 -199
rect 57 -203 63 -199
rect 73 -203 79 -199
rect 89 -203 95 -199
rect 42 -222 46 -218
rect 58 -222 62 -218
rect 74 -222 78 -218
rect 90 -222 94 -218
rect 315 -219 319 -197
rect 41 -235 47 -231
rect 57 -235 63 -231
rect 73 -235 79 -231
rect 89 -235 95 -231
rect 347 -154 351 -133
rect 347 -193 351 -169
rect 331 -219 335 -197
<< m2contact >>
rect 16 12 20 16
rect 34 12 38 16
rect 8 8 12 12
rect 42 12 46 16
rect 50 12 54 16
rect 58 12 62 16
rect 66 12 70 16
rect 74 12 78 16
rect 82 12 86 16
rect 90 12 94 16
rect 26 1 30 5
rect 98 -6 102 -2
rect 120 0 124 4
rect 98 -22 102 -18
rect 120 -16 124 -12
rect 98 -38 102 -34
rect 120 -32 124 -28
rect 26 -53 30 -49
rect 8 -60 12 -56
rect 1 -173 5 -169
rect 35 -65 39 -61
rect 43 -65 47 -61
rect 51 -65 55 -61
rect 59 -65 63 -61
rect 67 -65 71 -61
rect 75 -65 79 -61
rect 83 -65 87 -61
rect 91 -65 95 -61
rect 100 -64 104 -60
rect 137 -56 141 -52
rect 154 -8 158 -4
rect 276 15 280 19
rect 176 0 180 4
rect 199 -1 203 3
rect 306 24 310 28
rect 298 16 302 20
rect 350 16 354 20
rect 306 6 310 10
rect 261 -5 265 -1
rect 301 -5 305 -1
rect 154 -24 158 -20
rect 176 -16 180 -12
rect 199 -9 203 -5
rect 229 -13 233 -9
rect 199 -17 203 -13
rect 301 -13 305 -9
rect 261 -21 265 -17
rect 301 -21 305 -17
rect 154 -40 158 -36
rect 176 -32 180 -28
rect 199 -25 203 -21
rect 229 -29 233 -25
rect 199 -33 203 -29
rect 301 -29 305 -25
rect 348 6 352 10
rect 360 -5 364 -1
rect 360 -13 364 -9
rect 261 -37 265 -33
rect 301 -37 305 -33
rect 111 -72 115 -68
rect 8 -195 12 -191
rect 1 -203 5 -199
rect 8 -227 12 -223
rect 16 -86 20 -82
rect 100 -86 104 -82
rect 35 -110 39 -106
rect 51 -110 55 -106
rect 67 -110 71 -106
rect 83 -110 87 -106
rect 25 -173 29 -169
rect 43 -146 47 -142
rect 59 -146 63 -142
rect 75 -146 79 -142
rect 91 -146 95 -142
rect 111 -173 115 -169
rect 33 -185 37 -181
rect 41 -185 45 -181
rect 49 -185 53 -181
rect 57 -185 61 -181
rect 65 -185 69 -181
rect 73 -185 77 -181
rect 81 -185 85 -181
rect 89 -185 93 -181
rect 25 -195 29 -191
rect 100 -196 104 -192
rect 25 -203 29 -199
rect 42 -210 46 -206
rect 58 -210 62 -206
rect 74 -210 78 -206
rect 90 -210 94 -206
rect 34 -217 38 -213
rect 50 -217 54 -213
rect 66 -217 70 -213
rect 82 -217 86 -213
rect 25 -227 29 -223
rect 100 -228 104 -224
rect 42 -244 46 -240
rect 58 -244 62 -240
rect 74 -244 78 -240
rect 90 -244 94 -240
rect 100 -258 104 -254
rect 34 -269 38 -265
rect 50 -269 54 -265
rect 66 -269 70 -265
rect 82 -269 86 -265
rect 119 -64 123 -60
rect 147 -64 151 -60
rect 161 -64 165 -60
rect 199 -41 203 -37
rect 229 -45 233 -41
rect 192 -72 196 -68
rect 301 -45 305 -41
rect 236 -72 240 -68
rect 276 -56 280 -52
rect 315 -54 319 -50
rect 360 -21 364 -17
rect 360 -29 364 -25
rect 360 -37 364 -33
rect 360 -45 364 -41
rect 331 -54 335 -50
rect 147 -86 151 -82
rect 283 -64 287 -60
rect 276 -78 280 -74
rect 268 -130 272 -126
rect 126 -196 130 -192
rect 126 -228 130 -224
rect 119 -258 123 -254
rect 276 -249 280 -245
rect 307 -78 311 -74
rect 315 -98 319 -94
rect 331 -98 335 -94
rect 307 -130 311 -126
rect 323 -166 327 -162
rect 339 -166 343 -162
rect 307 -173 311 -169
rect 315 -228 319 -224
rect 331 -228 335 -224
rect 307 -249 311 -245
<< psubstratepcontact >>
rect 29 26 97 30
rect 348 0 352 4
rect 283 -5 287 -1
rect 348 -16 352 -12
rect 283 -21 287 -17
rect 348 -32 352 -28
rect 283 -37 287 -33
rect 348 -48 352 -44
rect 283 -56 291 -52
rect 315 -61 319 -57
rect 331 -61 335 -57
rect 35 -86 39 -82
rect 51 -86 55 -82
rect 67 -86 71 -82
rect 347 -61 351 -57
rect 83 -86 87 -82
rect 32 -251 36 -247
rect 48 -251 52 -247
rect 64 -251 68 -247
rect 80 -251 84 -247
rect 96 -251 100 -247
rect 315 -265 319 -261
rect 331 -265 335 -261
rect 347 -265 351 -261
<< nsubstratencontact >>
rect 313 29 345 33
rect 106 8 110 12
rect 0 -48 4 0
rect 192 8 196 12
rect 106 -8 110 -4
rect 192 -8 196 -4
rect 231 -5 235 -1
rect 106 -24 110 -20
rect 192 -24 196 -20
rect 231 -21 235 -17
rect 106 -40 110 -36
rect 192 -40 196 -36
rect 231 -37 235 -33
rect 35 -146 39 -142
rect 51 -146 55 -142
rect 67 -146 71 -142
rect 83 -146 87 -142
rect 315 -159 319 -155
rect 331 -159 335 -155
rect 32 -203 36 -199
rect 48 -203 52 -199
rect 64 -203 68 -199
rect 80 -203 84 -199
rect 96 -203 100 -199
rect 32 -235 36 -231
rect 48 -235 52 -231
rect 64 -235 68 -231
rect 80 -235 84 -231
rect 96 -235 100 -231
rect 347 -159 351 -155
<< labels >>
rlabel metal2 42 -246 45 -246 1 x
rlabel metal2 58 -246 61 -246 1 InSt0*
rlabel metal2 74 -246 77 -246 1 InSt1*
rlabel metal2 90 -246 93 -246 1 InSt2*
rlabel metal1 268 -264 271 -264 1 p1-
rlabel metal1 276 -264 279 -264 1 p1
rlabel metal1 127 -267 130 -267 1 p2-
rlabel metal1 119 -267 122 -267 1 p2
rlabel metal1 107 -267 115 -267 1 Vdd!
rlabel metal1 283 -264 291 -264 1 GND!
rlabel metal1 315 -222 318 -222 1 OutSt2*
rlabel metal2 323 -222 326 -222 1 OutSt1*
rlabel metal1 331 -222 334 -222 1 OutSt0*
rlabel metal2 339 -222 342 -222 1 z
<< end >>
