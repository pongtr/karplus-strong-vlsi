magic
tech scmos
timestamp 1512534937
use sreg_left_control  sreg_left_control_0
timestamp 1512534937
transform 1 0 -99 0 1 1181
box 4 -1178 99 65
use sreg  sreg_0
array 0 0 27 0 9 124
timestamp 1512338440
transform 1 0 9 0 1 100
box -9 -97 18 27
use sreg_01_right  sreg_01_right_0
array 0 0 19 0 9 124
timestamp 1512383252
transform 1 0 27 0 1 36
box -6 -33 15 95
<< end >>
