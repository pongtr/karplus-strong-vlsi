magic
tech scmos
timestamp 1512539734
<< polysilicon >>
rect -74 1238 -72 1240
rect -66 1238 -64 1240
rect -58 1238 -56 1240
rect -58 1170 -56 1172
<< metal1 >>
rect -95 1233 -93 1236
<< metal2 >>
rect -95 1222 -93 1226
rect -95 1127 -92 1131
rect 119 1127 121 1131
rect -95 1003 -93 1007
rect 119 1003 121 1007
rect -95 879 -93 883
rect 119 879 121 883
rect -95 755 -93 759
rect 119 755 121 759
rect -95 631 -93 635
rect 119 631 121 635
rect -95 507 -93 511
rect 119 507 121 511
rect -95 383 -93 387
rect 119 383 121 387
rect -95 259 -93 263
rect 119 259 121 263
rect -95 135 -93 139
rect 119 135 121 139
rect -95 11 -93 15
rect 119 11 121 15
use sreg_left_control  sreg_left_control_0
timestamp 1512534937
transform 1 0 -99 0 1 1181
box 4 -1178 99 65
use sreg_10b  sreg_10b_0
array 0 1 56 0 0 1248
timestamp 1512379799
transform 1 0 0 0 1 3
box 0 -3 56 1245
use sreg_right  sreg_right_0
timestamp 1512379879
transform 1 0 123 0 1 2
box -11 2 -2 1155
<< labels >>
rlabel metal1 -94 1233 -94 1236 3 Vdd!
rlabel metal2 -94 1222 -94 1226 3 GND!
rlabel polysilicon -74 1239 -72 1239 1 en
rlabel polysilicon -66 1239 -64 1239 1 bp
rlabel polysilicon -58 1239 -56 1239 1 phi0
rlabel polysilicon -58 1171 -56 1171 1 phi1
rlabel metal2 -94 1127 -94 1131 3 in9
rlabel metal2 120 1127 120 1131 7 out9
rlabel metal2 -94 1003 -94 1007 3 in8
rlabel metal2 -94 879 -94 883 3 in7
rlabel metal2 -94 755 -94 759 3 in6
rlabel metal2 -94 631 -94 635 3 in5
rlabel metal2 -94 507 -94 511 3 in4
rlabel metal2 -94 11 -94 15 3 in0
rlabel metal2 -94 135 -94 139 3 in1
rlabel metal2 -94 259 -94 263 3 in2
rlabel metal2 -94 383 -94 387 3 in3
rlabel metal2 120 1003 120 1007 7 out8
rlabel metal2 120 879 120 883 7 out7
rlabel metal2 120 755 120 759 7 out6
rlabel metal2 120 631 120 635 7 out5
rlabel metal2 120 11 120 15 7 out0
rlabel metal2 120 135 120 139 7 out1
rlabel metal2 120 259 120 263 7 out2
rlabel metal2 120 383 120 387 7 out3
rlabel metal2 120 507 120 511 7 out4
<< end >>
