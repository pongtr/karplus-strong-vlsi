magic
tech scmos
timestamp 1012241868
<< psubstratepdiff >>
rect 394 58 774 62
rect 394 54 541 58
rect 545 54 546 58
rect 550 54 551 58
rect 555 54 556 58
rect 560 54 570 58
rect 574 54 575 58
rect 579 54 580 58
rect 584 54 585 58
rect 589 54 599 58
rect 603 54 604 58
rect 608 54 609 58
rect 613 54 614 58
rect 618 54 628 58
rect 632 54 633 58
rect 637 54 638 58
rect 642 54 643 58
rect 647 54 657 58
rect 661 54 662 58
rect 666 54 667 58
rect 671 54 672 58
rect 676 54 774 58
rect 394 48 774 54
rect 394 44 541 48
rect 545 44 546 48
rect 550 44 551 48
rect 555 44 556 48
rect 560 44 570 48
rect 574 44 575 48
rect 579 44 580 48
rect 584 44 585 48
rect 589 44 599 48
rect 603 44 604 48
rect 608 44 609 48
rect 613 44 614 48
rect 618 44 628 48
rect 632 44 633 48
rect 637 44 638 48
rect 642 44 643 48
rect 647 44 657 48
rect 661 44 662 48
rect 666 44 667 48
rect 671 44 672 48
rect 676 44 774 48
rect 394 38 774 44
rect 394 34 541 38
rect 545 34 546 38
rect 550 34 551 38
rect 555 34 556 38
rect 560 34 570 38
rect 574 34 575 38
rect 579 34 580 38
rect 584 34 585 38
rect 589 34 599 38
rect 603 34 604 38
rect 608 34 609 38
rect 613 34 614 38
rect 618 34 628 38
rect 632 34 633 38
rect 637 34 638 38
rect 642 34 643 38
rect 647 34 657 38
rect 661 34 662 38
rect 666 34 667 38
rect 671 34 672 38
rect 676 34 774 38
rect 394 28 774 34
rect 394 24 541 28
rect 545 24 546 28
rect 550 24 551 28
rect 555 24 556 28
rect 560 24 570 28
rect 574 24 575 28
rect 579 24 580 28
rect 584 24 585 28
rect 589 24 599 28
rect 603 24 604 28
rect 608 24 609 28
rect 613 24 614 28
rect 618 24 628 28
rect 632 24 633 28
rect 637 24 638 28
rect 642 24 643 28
rect 647 24 657 28
rect 661 24 662 28
rect 666 24 667 28
rect 671 24 672 28
rect 676 24 774 28
rect 394 22 774 24
rect 394 -40 434 22
rect 394 -44 398 -40
rect 402 -44 408 -40
rect 412 -44 418 -40
rect 422 -44 428 -40
rect 432 -44 434 -40
rect 394 -45 434 -44
rect 394 -49 398 -45
rect 402 -49 408 -45
rect 412 -49 418 -45
rect 422 -49 428 -45
rect 432 -49 434 -45
rect 394 -50 434 -49
rect 394 -54 398 -50
rect 402 -54 408 -50
rect 412 -54 418 -50
rect 422 -54 428 -50
rect 432 -54 434 -50
rect 394 -55 434 -54
rect 394 -59 398 -55
rect 402 -59 408 -55
rect 412 -59 418 -55
rect 422 -59 428 -55
rect 432 -59 434 -55
rect 394 -66 434 -59
rect 394 -70 398 -66
rect 402 -70 408 -66
rect 412 -70 418 -66
rect 422 -70 428 -66
rect 432 -70 434 -66
rect 394 -71 434 -70
rect 394 -75 398 -71
rect 402 -75 408 -71
rect 412 -75 418 -71
rect 422 -75 428 -71
rect 432 -75 434 -71
rect 394 -76 434 -75
rect 394 -80 398 -76
rect 402 -80 408 -76
rect 412 -80 418 -76
rect 422 -80 428 -76
rect 432 -80 434 -76
rect 394 -81 434 -80
rect 394 -85 398 -81
rect 402 -85 408 -81
rect 412 -85 418 -81
rect 422 -85 428 -81
rect 432 -85 434 -81
rect 394 -92 434 -85
rect 394 -96 398 -92
rect 402 -96 408 -92
rect 412 -96 418 -92
rect 422 -96 428 -92
rect 432 -96 434 -92
rect 394 -97 434 -96
rect 394 -101 398 -97
rect 402 -101 408 -97
rect 412 -101 418 -97
rect 422 -101 428 -97
rect 432 -101 434 -97
rect 394 -102 434 -101
rect 394 -106 398 -102
rect 402 -106 408 -102
rect 412 -106 418 -102
rect 422 -106 428 -102
rect 432 -106 434 -102
rect 394 -107 434 -106
rect 394 -111 398 -107
rect 402 -111 408 -107
rect 412 -111 418 -107
rect 422 -111 428 -107
rect 432 -111 434 -107
rect 394 -118 434 -111
rect 394 -122 398 -118
rect 402 -122 408 -118
rect 412 -122 418 -118
rect 422 -122 428 -118
rect 432 -122 434 -118
rect 394 -123 434 -122
rect 394 -127 398 -123
rect 402 -127 408 -123
rect 412 -127 418 -123
rect 422 -127 428 -123
rect 432 -127 434 -123
rect 394 -128 434 -127
rect 394 -132 398 -128
rect 402 -132 408 -128
rect 412 -132 418 -128
rect 422 -132 428 -128
rect 432 -132 434 -128
rect 394 -133 434 -132
rect 394 -137 398 -133
rect 402 -137 408 -133
rect 412 -137 418 -133
rect 422 -137 428 -133
rect 432 -137 434 -133
rect 394 -144 434 -137
rect 394 -148 398 -144
rect 402 -148 408 -144
rect 412 -148 418 -144
rect 422 -148 428 -144
rect 432 -148 434 -144
rect 394 -149 434 -148
rect 394 -153 398 -149
rect 402 -153 408 -149
rect 412 -153 418 -149
rect 422 -153 428 -149
rect 432 -153 434 -149
rect 394 -154 434 -153
rect 394 -158 398 -154
rect 402 -158 408 -154
rect 412 -158 418 -154
rect 422 -158 428 -154
rect 432 -158 434 -154
rect 394 -159 434 -158
rect 394 -163 398 -159
rect 402 -163 408 -159
rect 412 -163 418 -159
rect 422 -163 428 -159
rect 432 -163 434 -159
rect 394 -331 434 -163
<< nsubstratendiff >>
rect 348 104 774 108
rect 348 100 541 104
rect 545 100 546 104
rect 550 100 551 104
rect 555 100 556 104
rect 560 100 570 104
rect 574 100 575 104
rect 579 100 580 104
rect 584 100 585 104
rect 589 100 599 104
rect 603 100 604 104
rect 608 100 609 104
rect 613 100 614 104
rect 618 100 628 104
rect 632 100 633 104
rect 637 100 638 104
rect 642 100 643 104
rect 647 100 657 104
rect 661 100 662 104
rect 666 100 667 104
rect 671 100 672 104
rect 676 100 774 104
rect 348 94 774 100
rect 348 90 541 94
rect 545 90 546 94
rect 550 90 551 94
rect 555 90 556 94
rect 560 90 570 94
rect 574 90 575 94
rect 579 90 580 94
rect 584 90 585 94
rect 589 90 599 94
rect 603 90 604 94
rect 608 90 609 94
rect 613 90 614 94
rect 618 90 628 94
rect 632 90 633 94
rect 637 90 638 94
rect 642 90 643 94
rect 647 90 657 94
rect 661 90 662 94
rect 666 90 667 94
rect 671 90 672 94
rect 676 90 774 94
rect 348 84 774 90
rect 348 80 541 84
rect 545 80 546 84
rect 550 80 551 84
rect 555 80 556 84
rect 560 80 570 84
rect 574 80 575 84
rect 579 80 580 84
rect 584 80 585 84
rect 589 80 599 84
rect 603 80 604 84
rect 608 80 609 84
rect 613 80 614 84
rect 618 80 628 84
rect 632 80 633 84
rect 637 80 638 84
rect 642 80 643 84
rect 647 80 657 84
rect 661 80 662 84
rect 666 80 667 84
rect 671 80 672 84
rect 676 80 774 84
rect 348 74 774 80
rect 348 70 541 74
rect 545 70 546 74
rect 550 70 551 74
rect 555 70 556 74
rect 560 70 570 74
rect 574 70 575 74
rect 579 70 580 74
rect 584 70 585 74
rect 589 70 599 74
rect 603 70 604 74
rect 608 70 609 74
rect 613 70 614 74
rect 618 70 628 74
rect 632 70 633 74
rect 637 70 638 74
rect 642 70 643 74
rect 647 70 657 74
rect 661 70 662 74
rect 666 70 667 74
rect 671 70 672 74
rect 676 70 774 74
rect 348 68 774 70
rect 348 -40 388 68
rect 348 -44 352 -40
rect 356 -44 362 -40
rect 366 -44 372 -40
rect 376 -44 382 -40
rect 386 -44 388 -40
rect 348 -45 388 -44
rect 348 -49 352 -45
rect 356 -49 362 -45
rect 366 -49 372 -45
rect 376 -49 382 -45
rect 386 -49 388 -45
rect 348 -50 388 -49
rect 348 -54 352 -50
rect 356 -54 362 -50
rect 366 -54 372 -50
rect 376 -54 382 -50
rect 386 -54 388 -50
rect 348 -55 388 -54
rect 348 -59 352 -55
rect 356 -59 362 -55
rect 366 -59 372 -55
rect 376 -59 382 -55
rect 386 -59 388 -55
rect 348 -66 388 -59
rect 348 -70 352 -66
rect 356 -70 362 -66
rect 366 -70 372 -66
rect 376 -70 382 -66
rect 386 -70 388 -66
rect 348 -71 388 -70
rect 348 -75 352 -71
rect 356 -75 362 -71
rect 366 -75 372 -71
rect 376 -75 382 -71
rect 386 -75 388 -71
rect 348 -76 388 -75
rect 348 -80 352 -76
rect 356 -80 362 -76
rect 366 -80 372 -76
rect 376 -80 382 -76
rect 386 -80 388 -76
rect 348 -81 388 -80
rect 348 -85 352 -81
rect 356 -85 362 -81
rect 366 -85 372 -81
rect 376 -85 382 -81
rect 386 -85 388 -81
rect 348 -92 388 -85
rect 348 -96 352 -92
rect 356 -96 362 -92
rect 366 -96 372 -92
rect 376 -96 382 -92
rect 386 -96 388 -92
rect 348 -97 388 -96
rect 348 -101 352 -97
rect 356 -101 362 -97
rect 366 -101 372 -97
rect 376 -101 382 -97
rect 386 -101 388 -97
rect 348 -102 388 -101
rect 348 -106 352 -102
rect 356 -106 362 -102
rect 366 -106 372 -102
rect 376 -106 382 -102
rect 386 -106 388 -102
rect 348 -107 388 -106
rect 348 -111 352 -107
rect 356 -111 362 -107
rect 366 -111 372 -107
rect 376 -111 382 -107
rect 386 -111 388 -107
rect 348 -118 388 -111
rect 348 -122 352 -118
rect 356 -122 362 -118
rect 366 -122 372 -118
rect 376 -122 382 -118
rect 386 -122 388 -118
rect 348 -123 388 -122
rect 348 -127 352 -123
rect 356 -127 362 -123
rect 366 -127 372 -123
rect 376 -127 382 -123
rect 386 -127 388 -123
rect 348 -128 388 -127
rect 348 -132 352 -128
rect 356 -132 362 -128
rect 366 -132 372 -128
rect 376 -132 382 -128
rect 386 -132 388 -128
rect 348 -133 388 -132
rect 348 -137 352 -133
rect 356 -137 362 -133
rect 366 -137 372 -133
rect 376 -137 382 -133
rect 386 -137 388 -133
rect 348 -144 388 -137
rect 348 -148 352 -144
rect 356 -148 362 -144
rect 366 -148 372 -144
rect 376 -148 382 -144
rect 386 -148 388 -144
rect 348 -149 388 -148
rect 348 -153 352 -149
rect 356 -153 362 -149
rect 366 -153 372 -149
rect 376 -153 382 -149
rect 386 -153 388 -149
rect 348 -154 388 -153
rect 348 -158 352 -154
rect 356 -158 362 -154
rect 366 -158 372 -154
rect 376 -158 382 -154
rect 386 -158 388 -154
rect 348 -159 388 -158
rect 348 -163 352 -159
rect 356 -163 362 -159
rect 366 -163 372 -159
rect 376 -163 382 -159
rect 386 -163 388 -159
rect 348 -331 388 -163
<< psubstratepcontact >>
rect 541 54 545 58
rect 546 54 550 58
rect 551 54 555 58
rect 556 54 560 58
rect 570 54 574 58
rect 575 54 579 58
rect 580 54 584 58
rect 585 54 589 58
rect 599 54 603 58
rect 604 54 608 58
rect 609 54 613 58
rect 614 54 618 58
rect 628 54 632 58
rect 633 54 637 58
rect 638 54 642 58
rect 643 54 647 58
rect 657 54 661 58
rect 662 54 666 58
rect 667 54 671 58
rect 672 54 676 58
rect 541 44 545 48
rect 546 44 550 48
rect 551 44 555 48
rect 556 44 560 48
rect 570 44 574 48
rect 575 44 579 48
rect 580 44 584 48
rect 585 44 589 48
rect 599 44 603 48
rect 604 44 608 48
rect 609 44 613 48
rect 614 44 618 48
rect 628 44 632 48
rect 633 44 637 48
rect 638 44 642 48
rect 643 44 647 48
rect 657 44 661 48
rect 662 44 666 48
rect 667 44 671 48
rect 672 44 676 48
rect 541 34 545 38
rect 546 34 550 38
rect 551 34 555 38
rect 556 34 560 38
rect 570 34 574 38
rect 575 34 579 38
rect 580 34 584 38
rect 585 34 589 38
rect 599 34 603 38
rect 604 34 608 38
rect 609 34 613 38
rect 614 34 618 38
rect 628 34 632 38
rect 633 34 637 38
rect 638 34 642 38
rect 643 34 647 38
rect 657 34 661 38
rect 662 34 666 38
rect 667 34 671 38
rect 672 34 676 38
rect 541 24 545 28
rect 546 24 550 28
rect 551 24 555 28
rect 556 24 560 28
rect 570 24 574 28
rect 575 24 579 28
rect 580 24 584 28
rect 585 24 589 28
rect 599 24 603 28
rect 604 24 608 28
rect 609 24 613 28
rect 614 24 618 28
rect 628 24 632 28
rect 633 24 637 28
rect 638 24 642 28
rect 643 24 647 28
rect 657 24 661 28
rect 662 24 666 28
rect 667 24 671 28
rect 672 24 676 28
rect 398 -44 402 -40
rect 408 -44 412 -40
rect 418 -44 422 -40
rect 428 -44 432 -40
rect 398 -49 402 -45
rect 408 -49 412 -45
rect 418 -49 422 -45
rect 428 -49 432 -45
rect 398 -54 402 -50
rect 408 -54 412 -50
rect 418 -54 422 -50
rect 428 -54 432 -50
rect 398 -59 402 -55
rect 408 -59 412 -55
rect 418 -59 422 -55
rect 428 -59 432 -55
rect 398 -70 402 -66
rect 408 -70 412 -66
rect 418 -70 422 -66
rect 428 -70 432 -66
rect 398 -75 402 -71
rect 408 -75 412 -71
rect 418 -75 422 -71
rect 428 -75 432 -71
rect 398 -80 402 -76
rect 408 -80 412 -76
rect 418 -80 422 -76
rect 428 -80 432 -76
rect 398 -85 402 -81
rect 408 -85 412 -81
rect 418 -85 422 -81
rect 428 -85 432 -81
rect 398 -96 402 -92
rect 408 -96 412 -92
rect 418 -96 422 -92
rect 428 -96 432 -92
rect 398 -101 402 -97
rect 408 -101 412 -97
rect 418 -101 422 -97
rect 428 -101 432 -97
rect 398 -106 402 -102
rect 408 -106 412 -102
rect 418 -106 422 -102
rect 428 -106 432 -102
rect 398 -111 402 -107
rect 408 -111 412 -107
rect 418 -111 422 -107
rect 428 -111 432 -107
rect 398 -122 402 -118
rect 408 -122 412 -118
rect 418 -122 422 -118
rect 428 -122 432 -118
rect 398 -127 402 -123
rect 408 -127 412 -123
rect 418 -127 422 -123
rect 428 -127 432 -123
rect 398 -132 402 -128
rect 408 -132 412 -128
rect 418 -132 422 -128
rect 428 -132 432 -128
rect 398 -137 402 -133
rect 408 -137 412 -133
rect 418 -137 422 -133
rect 428 -137 432 -133
rect 398 -148 402 -144
rect 408 -148 412 -144
rect 418 -148 422 -144
rect 428 -148 432 -144
rect 398 -153 402 -149
rect 408 -153 412 -149
rect 418 -153 422 -149
rect 428 -153 432 -149
rect 398 -158 402 -154
rect 408 -158 412 -154
rect 418 -158 422 -154
rect 428 -158 432 -154
rect 398 -163 402 -159
rect 408 -163 412 -159
rect 418 -163 422 -159
rect 428 -163 432 -159
<< nsubstratencontact >>
rect 541 100 545 104
rect 546 100 550 104
rect 551 100 555 104
rect 556 100 560 104
rect 570 100 574 104
rect 575 100 579 104
rect 580 100 584 104
rect 585 100 589 104
rect 599 100 603 104
rect 604 100 608 104
rect 609 100 613 104
rect 614 100 618 104
rect 628 100 632 104
rect 633 100 637 104
rect 638 100 642 104
rect 643 100 647 104
rect 657 100 661 104
rect 662 100 666 104
rect 667 100 671 104
rect 672 100 676 104
rect 541 90 545 94
rect 546 90 550 94
rect 551 90 555 94
rect 556 90 560 94
rect 570 90 574 94
rect 575 90 579 94
rect 580 90 584 94
rect 585 90 589 94
rect 599 90 603 94
rect 604 90 608 94
rect 609 90 613 94
rect 614 90 618 94
rect 628 90 632 94
rect 633 90 637 94
rect 638 90 642 94
rect 643 90 647 94
rect 657 90 661 94
rect 662 90 666 94
rect 667 90 671 94
rect 672 90 676 94
rect 541 80 545 84
rect 546 80 550 84
rect 551 80 555 84
rect 556 80 560 84
rect 570 80 574 84
rect 575 80 579 84
rect 580 80 584 84
rect 585 80 589 84
rect 599 80 603 84
rect 604 80 608 84
rect 609 80 613 84
rect 614 80 618 84
rect 628 80 632 84
rect 633 80 637 84
rect 638 80 642 84
rect 643 80 647 84
rect 657 80 661 84
rect 662 80 666 84
rect 667 80 671 84
rect 672 80 676 84
rect 541 70 545 74
rect 546 70 550 74
rect 551 70 555 74
rect 556 70 560 74
rect 570 70 574 74
rect 575 70 579 74
rect 580 70 584 74
rect 585 70 589 74
rect 599 70 603 74
rect 604 70 608 74
rect 609 70 613 74
rect 614 70 618 74
rect 628 70 632 74
rect 633 70 637 74
rect 638 70 642 74
rect 643 70 647 74
rect 657 70 661 74
rect 662 70 666 74
rect 667 70 671 74
rect 672 70 676 74
rect 352 -44 356 -40
rect 362 -44 366 -40
rect 372 -44 376 -40
rect 382 -44 386 -40
rect 352 -49 356 -45
rect 362 -49 366 -45
rect 372 -49 376 -45
rect 382 -49 386 -45
rect 352 -54 356 -50
rect 362 -54 366 -50
rect 372 -54 376 -50
rect 382 -54 386 -50
rect 352 -59 356 -55
rect 362 -59 366 -55
rect 372 -59 376 -55
rect 382 -59 386 -55
rect 352 -70 356 -66
rect 362 -70 366 -66
rect 372 -70 376 -66
rect 382 -70 386 -66
rect 352 -75 356 -71
rect 362 -75 366 -71
rect 372 -75 376 -71
rect 382 -75 386 -71
rect 352 -80 356 -76
rect 362 -80 366 -76
rect 372 -80 376 -76
rect 382 -80 386 -76
rect 352 -85 356 -81
rect 362 -85 366 -81
rect 372 -85 376 -81
rect 382 -85 386 -81
rect 352 -96 356 -92
rect 362 -96 366 -92
rect 372 -96 376 -92
rect 382 -96 386 -92
rect 352 -101 356 -97
rect 362 -101 366 -97
rect 372 -101 376 -97
rect 382 -101 386 -97
rect 352 -106 356 -102
rect 362 -106 366 -102
rect 372 -106 376 -102
rect 382 -106 386 -102
rect 352 -111 356 -107
rect 362 -111 366 -107
rect 372 -111 376 -107
rect 382 -111 386 -107
rect 352 -122 356 -118
rect 362 -122 366 -118
rect 372 -122 376 -118
rect 382 -122 386 -118
rect 352 -127 356 -123
rect 362 -127 366 -123
rect 372 -127 376 -123
rect 382 -127 386 -123
rect 352 -132 356 -128
rect 362 -132 366 -128
rect 372 -132 376 -128
rect 382 -132 386 -128
rect 352 -137 356 -133
rect 362 -137 366 -133
rect 372 -137 376 -133
rect 382 -137 386 -133
rect 352 -148 356 -144
rect 362 -148 366 -144
rect 372 -148 376 -144
rect 382 -148 386 -144
rect 352 -153 356 -149
rect 362 -153 366 -149
rect 372 -153 376 -149
rect 382 -153 386 -149
rect 352 -158 356 -154
rect 362 -158 366 -154
rect 372 -158 376 -154
rect 382 -158 386 -154
rect 352 -163 356 -159
rect 362 -163 366 -159
rect 372 -163 376 -159
rect 382 -163 386 -159
<< polysilicon >>
rect -143 124 763 618
rect -143 -314 332 124
<< metal1 >>
rect -143 124 763 618
rect -143 -314 332 124
rect 545 100 546 104
rect 550 100 551 104
rect 555 100 556 104
rect 541 99 560 100
rect 545 95 546 99
rect 550 95 551 99
rect 555 95 556 99
rect 541 94 560 95
rect 545 90 546 94
rect 550 90 551 94
rect 555 90 556 94
rect 541 89 560 90
rect 545 85 546 89
rect 550 85 551 89
rect 555 85 556 89
rect 541 84 560 85
rect 545 80 546 84
rect 550 80 551 84
rect 555 80 556 84
rect 541 79 560 80
rect 545 75 546 79
rect 550 75 551 79
rect 555 75 556 79
rect 541 74 560 75
rect 545 70 546 74
rect 550 70 551 74
rect 555 70 556 74
rect 574 100 575 104
rect 579 100 580 104
rect 584 100 585 104
rect 570 99 589 100
rect 574 95 575 99
rect 579 95 580 99
rect 584 95 585 99
rect 570 94 589 95
rect 574 90 575 94
rect 579 90 580 94
rect 584 90 585 94
rect 570 89 589 90
rect 574 85 575 89
rect 579 85 580 89
rect 584 85 585 89
rect 570 84 589 85
rect 574 80 575 84
rect 579 80 580 84
rect 584 80 585 84
rect 570 79 589 80
rect 574 75 575 79
rect 579 75 580 79
rect 584 75 585 79
rect 570 74 589 75
rect 574 70 575 74
rect 579 70 580 74
rect 584 70 585 74
rect 603 100 604 104
rect 608 100 609 104
rect 613 100 614 104
rect 599 99 618 100
rect 603 95 604 99
rect 608 95 609 99
rect 613 95 614 99
rect 599 94 618 95
rect 603 90 604 94
rect 608 90 609 94
rect 613 90 614 94
rect 599 89 618 90
rect 603 85 604 89
rect 608 85 609 89
rect 613 85 614 89
rect 599 84 618 85
rect 603 80 604 84
rect 608 80 609 84
rect 613 80 614 84
rect 599 79 618 80
rect 603 75 604 79
rect 608 75 609 79
rect 613 75 614 79
rect 599 74 618 75
rect 603 70 604 74
rect 608 70 609 74
rect 613 70 614 74
rect 632 100 633 104
rect 637 100 638 104
rect 642 100 643 104
rect 628 99 647 100
rect 632 95 633 99
rect 637 95 638 99
rect 642 95 643 99
rect 628 94 647 95
rect 632 90 633 94
rect 637 90 638 94
rect 642 90 643 94
rect 628 89 647 90
rect 632 85 633 89
rect 637 85 638 89
rect 642 85 643 89
rect 628 84 647 85
rect 632 80 633 84
rect 637 80 638 84
rect 642 80 643 84
rect 628 79 647 80
rect 632 75 633 79
rect 637 75 638 79
rect 642 75 643 79
rect 628 74 647 75
rect 632 70 633 74
rect 637 70 638 74
rect 642 70 643 74
rect 661 100 662 104
rect 666 100 667 104
rect 671 100 672 104
rect 657 99 676 100
rect 661 95 662 99
rect 666 95 667 99
rect 671 95 672 99
rect 657 94 676 95
rect 661 90 662 94
rect 666 90 667 94
rect 671 90 672 94
rect 657 89 676 90
rect 661 85 662 89
rect 666 85 667 89
rect 671 85 672 89
rect 657 84 676 85
rect 661 80 662 84
rect 666 80 667 84
rect 671 80 672 84
rect 657 79 676 80
rect 661 75 662 79
rect 666 75 667 79
rect 671 75 672 79
rect 657 74 676 75
rect 661 70 662 74
rect 666 70 667 74
rect 671 70 672 74
rect 545 54 546 58
rect 550 54 551 58
rect 555 54 556 58
rect 541 53 560 54
rect 545 49 546 53
rect 550 49 551 53
rect 555 49 556 53
rect 541 48 560 49
rect 545 44 546 48
rect 550 44 551 48
rect 555 44 556 48
rect 541 43 560 44
rect 545 39 546 43
rect 550 39 551 43
rect 555 39 556 43
rect 541 38 560 39
rect 545 34 546 38
rect 550 34 551 38
rect 555 34 556 38
rect 541 33 560 34
rect 545 29 546 33
rect 550 29 551 33
rect 555 29 556 33
rect 541 28 560 29
rect 545 24 546 28
rect 550 24 551 28
rect 555 24 556 28
rect 574 54 575 58
rect 579 54 580 58
rect 584 54 585 58
rect 570 53 589 54
rect 574 49 575 53
rect 579 49 580 53
rect 584 49 585 53
rect 570 48 589 49
rect 574 44 575 48
rect 579 44 580 48
rect 584 44 585 48
rect 570 43 589 44
rect 574 39 575 43
rect 579 39 580 43
rect 584 39 585 43
rect 570 38 589 39
rect 574 34 575 38
rect 579 34 580 38
rect 584 34 585 38
rect 570 33 589 34
rect 574 29 575 33
rect 579 29 580 33
rect 584 29 585 33
rect 570 28 589 29
rect 574 24 575 28
rect 579 24 580 28
rect 584 24 585 28
rect 603 54 604 58
rect 608 54 609 58
rect 613 54 614 58
rect 599 53 618 54
rect 603 49 604 53
rect 608 49 609 53
rect 613 49 614 53
rect 599 48 618 49
rect 603 44 604 48
rect 608 44 609 48
rect 613 44 614 48
rect 599 43 618 44
rect 603 39 604 43
rect 608 39 609 43
rect 613 39 614 43
rect 599 38 618 39
rect 603 34 604 38
rect 608 34 609 38
rect 613 34 614 38
rect 599 33 618 34
rect 603 29 604 33
rect 608 29 609 33
rect 613 29 614 33
rect 599 28 618 29
rect 603 24 604 28
rect 608 24 609 28
rect 613 24 614 28
rect 632 54 633 58
rect 637 54 638 58
rect 642 54 643 58
rect 628 53 647 54
rect 632 49 633 53
rect 637 49 638 53
rect 642 49 643 53
rect 628 48 647 49
rect 632 44 633 48
rect 637 44 638 48
rect 642 44 643 48
rect 628 43 647 44
rect 632 39 633 43
rect 637 39 638 43
rect 642 39 643 43
rect 628 38 647 39
rect 632 34 633 38
rect 637 34 638 38
rect 642 34 643 38
rect 628 33 647 34
rect 632 29 633 33
rect 637 29 638 33
rect 642 29 643 33
rect 628 28 647 29
rect 632 24 633 28
rect 637 24 638 28
rect 642 24 643 28
rect 661 54 662 58
rect 666 54 667 58
rect 671 54 672 58
rect 657 53 676 54
rect 661 49 662 53
rect 666 49 667 53
rect 671 49 672 53
rect 657 48 676 49
rect 661 44 662 48
rect 666 44 667 48
rect 671 44 672 48
rect 657 43 676 44
rect 661 39 662 43
rect 666 39 667 43
rect 671 39 672 43
rect 657 38 676 39
rect 661 34 662 38
rect 666 34 667 38
rect 671 34 672 38
rect 657 33 676 34
rect 661 29 662 33
rect 666 29 667 33
rect 671 29 672 33
rect 657 28 676 29
rect 661 24 662 28
rect 666 24 667 28
rect 671 24 672 28
rect 356 -44 357 -40
rect 361 -44 362 -40
rect 366 -44 367 -40
rect 371 -44 372 -40
rect 376 -44 377 -40
rect 381 -44 382 -40
rect 352 -45 386 -44
rect 356 -49 357 -45
rect 361 -49 362 -45
rect 366 -49 367 -45
rect 371 -49 372 -45
rect 376 -49 377 -45
rect 381 -49 382 -45
rect 352 -50 386 -49
rect 356 -54 357 -50
rect 361 -54 362 -50
rect 366 -54 367 -50
rect 371 -54 372 -50
rect 376 -54 377 -50
rect 381 -54 382 -50
rect 352 -55 386 -54
rect 356 -59 357 -55
rect 361 -59 362 -55
rect 366 -59 367 -55
rect 371 -59 372 -55
rect 376 -59 377 -55
rect 381 -59 382 -55
rect 402 -44 403 -40
rect 407 -44 408 -40
rect 412 -44 413 -40
rect 417 -44 418 -40
rect 422 -44 423 -40
rect 427 -44 428 -40
rect 398 -45 432 -44
rect 402 -49 403 -45
rect 407 -49 408 -45
rect 412 -49 413 -45
rect 417 -49 418 -45
rect 422 -49 423 -45
rect 427 -49 428 -45
rect 398 -50 432 -49
rect 402 -54 403 -50
rect 407 -54 408 -50
rect 412 -54 413 -50
rect 417 -54 418 -50
rect 422 -54 423 -50
rect 427 -54 428 -50
rect 398 -55 432 -54
rect 402 -59 403 -55
rect 407 -59 408 -55
rect 412 -59 413 -55
rect 417 -59 418 -55
rect 422 -59 423 -55
rect 427 -59 428 -55
rect 356 -70 357 -66
rect 361 -70 362 -66
rect 366 -70 367 -66
rect 371 -70 372 -66
rect 376 -70 377 -66
rect 381 -70 382 -66
rect 352 -71 386 -70
rect 356 -75 357 -71
rect 361 -75 362 -71
rect 366 -75 367 -71
rect 371 -75 372 -71
rect 376 -75 377 -71
rect 381 -75 382 -71
rect 352 -76 386 -75
rect 356 -80 357 -76
rect 361 -80 362 -76
rect 366 -80 367 -76
rect 371 -80 372 -76
rect 376 -80 377 -76
rect 381 -80 382 -76
rect 352 -81 386 -80
rect 356 -85 357 -81
rect 361 -85 362 -81
rect 366 -85 367 -81
rect 371 -85 372 -81
rect 376 -85 377 -81
rect 381 -85 382 -81
rect 402 -70 403 -66
rect 407 -70 408 -66
rect 412 -70 413 -66
rect 417 -70 418 -66
rect 422 -70 423 -66
rect 427 -70 428 -66
rect 398 -71 432 -70
rect 402 -75 403 -71
rect 407 -75 408 -71
rect 412 -75 413 -71
rect 417 -75 418 -71
rect 422 -75 423 -71
rect 427 -75 428 -71
rect 398 -76 432 -75
rect 402 -80 403 -76
rect 407 -80 408 -76
rect 412 -80 413 -76
rect 417 -80 418 -76
rect 422 -80 423 -76
rect 427 -80 428 -76
rect 398 -81 432 -80
rect 402 -85 403 -81
rect 407 -85 408 -81
rect 412 -85 413 -81
rect 417 -85 418 -81
rect 422 -85 423 -81
rect 427 -85 428 -81
rect 356 -96 357 -92
rect 361 -96 362 -92
rect 366 -96 367 -92
rect 371 -96 372 -92
rect 376 -96 377 -92
rect 381 -96 382 -92
rect 352 -97 386 -96
rect 356 -101 357 -97
rect 361 -101 362 -97
rect 366 -101 367 -97
rect 371 -101 372 -97
rect 376 -101 377 -97
rect 381 -101 382 -97
rect 352 -102 386 -101
rect 356 -106 357 -102
rect 361 -106 362 -102
rect 366 -106 367 -102
rect 371 -106 372 -102
rect 376 -106 377 -102
rect 381 -106 382 -102
rect 352 -107 386 -106
rect 356 -111 357 -107
rect 361 -111 362 -107
rect 366 -111 367 -107
rect 371 -111 372 -107
rect 376 -111 377 -107
rect 381 -111 382 -107
rect 402 -96 403 -92
rect 407 -96 408 -92
rect 412 -96 413 -92
rect 417 -96 418 -92
rect 422 -96 423 -92
rect 427 -96 428 -92
rect 398 -97 432 -96
rect 402 -101 403 -97
rect 407 -101 408 -97
rect 412 -101 413 -97
rect 417 -101 418 -97
rect 422 -101 423 -97
rect 427 -101 428 -97
rect 398 -102 432 -101
rect 402 -106 403 -102
rect 407 -106 408 -102
rect 412 -106 413 -102
rect 417 -106 418 -102
rect 422 -106 423 -102
rect 427 -106 428 -102
rect 398 -107 432 -106
rect 402 -111 403 -107
rect 407 -111 408 -107
rect 412 -111 413 -107
rect 417 -111 418 -107
rect 422 -111 423 -107
rect 427 -111 428 -107
rect 356 -122 357 -118
rect 361 -122 362 -118
rect 366 -122 367 -118
rect 371 -122 372 -118
rect 376 -122 377 -118
rect 381 -122 382 -118
rect 352 -123 386 -122
rect 356 -127 357 -123
rect 361 -127 362 -123
rect 366 -127 367 -123
rect 371 -127 372 -123
rect 376 -127 377 -123
rect 381 -127 382 -123
rect 352 -128 386 -127
rect 356 -132 357 -128
rect 361 -132 362 -128
rect 366 -132 367 -128
rect 371 -132 372 -128
rect 376 -132 377 -128
rect 381 -132 382 -128
rect 352 -133 386 -132
rect 356 -137 357 -133
rect 361 -137 362 -133
rect 366 -137 367 -133
rect 371 -137 372 -133
rect 376 -137 377 -133
rect 381 -137 382 -133
rect 402 -122 403 -118
rect 407 -122 408 -118
rect 412 -122 413 -118
rect 417 -122 418 -118
rect 422 -122 423 -118
rect 427 -122 428 -118
rect 398 -123 432 -122
rect 402 -127 403 -123
rect 407 -127 408 -123
rect 412 -127 413 -123
rect 417 -127 418 -123
rect 422 -127 423 -123
rect 427 -127 428 -123
rect 398 -128 432 -127
rect 402 -132 403 -128
rect 407 -132 408 -128
rect 412 -132 413 -128
rect 417 -132 418 -128
rect 422 -132 423 -128
rect 427 -132 428 -128
rect 398 -133 432 -132
rect 402 -137 403 -133
rect 407 -137 408 -133
rect 412 -137 413 -133
rect 417 -137 418 -133
rect 422 -137 423 -133
rect 427 -137 428 -133
rect 356 -148 357 -144
rect 361 -148 362 -144
rect 366 -148 367 -144
rect 371 -148 372 -144
rect 376 -148 377 -144
rect 381 -148 382 -144
rect 352 -149 386 -148
rect 356 -153 357 -149
rect 361 -153 362 -149
rect 366 -153 367 -149
rect 371 -153 372 -149
rect 376 -153 377 -149
rect 381 -153 382 -149
rect 352 -154 386 -153
rect 356 -158 357 -154
rect 361 -158 362 -154
rect 366 -158 367 -154
rect 371 -158 372 -154
rect 376 -158 377 -154
rect 381 -158 382 -154
rect 352 -159 386 -158
rect 356 -163 357 -159
rect 361 -163 362 -159
rect 366 -163 367 -159
rect 371 -163 372 -159
rect 376 -163 377 -159
rect 381 -163 382 -159
rect 402 -148 403 -144
rect 407 -148 408 -144
rect 412 -148 413 -144
rect 417 -148 418 -144
rect 422 -148 423 -144
rect 427 -148 428 -144
rect 398 -149 432 -148
rect 402 -153 403 -149
rect 407 -153 408 -149
rect 412 -153 413 -149
rect 417 -153 418 -149
rect 422 -153 423 -149
rect 427 -153 428 -149
rect 398 -154 432 -153
rect 402 -158 403 -154
rect 407 -158 408 -154
rect 412 -158 413 -154
rect 417 -158 418 -154
rect 422 -158 423 -154
rect 427 -158 428 -154
rect 398 -159 432 -158
rect 402 -163 403 -159
rect 407 -163 408 -159
rect 412 -163 413 -159
rect 417 -163 418 -159
rect 422 -163 423 -159
rect 427 -163 428 -159
<< m2contact >>
rect 541 95 545 99
rect 546 95 550 99
rect 551 95 555 99
rect 556 95 560 99
rect 541 85 545 89
rect 546 85 550 89
rect 551 85 555 89
rect 556 85 560 89
rect 541 75 545 79
rect 546 75 550 79
rect 551 75 555 79
rect 556 75 560 79
rect 570 95 574 99
rect 575 95 579 99
rect 580 95 584 99
rect 585 95 589 99
rect 570 85 574 89
rect 575 85 579 89
rect 580 85 584 89
rect 585 85 589 89
rect 570 75 574 79
rect 575 75 579 79
rect 580 75 584 79
rect 585 75 589 79
rect 599 95 603 99
rect 604 95 608 99
rect 609 95 613 99
rect 614 95 618 99
rect 599 85 603 89
rect 604 85 608 89
rect 609 85 613 89
rect 614 85 618 89
rect 599 75 603 79
rect 604 75 608 79
rect 609 75 613 79
rect 614 75 618 79
rect 628 95 632 99
rect 633 95 637 99
rect 638 95 642 99
rect 643 95 647 99
rect 628 85 632 89
rect 633 85 637 89
rect 638 85 642 89
rect 643 85 647 89
rect 628 75 632 79
rect 633 75 637 79
rect 638 75 642 79
rect 643 75 647 79
rect 657 95 661 99
rect 662 95 666 99
rect 667 95 671 99
rect 672 95 676 99
rect 657 85 661 89
rect 662 85 666 89
rect 667 85 671 89
rect 672 85 676 89
rect 657 75 661 79
rect 662 75 666 79
rect 667 75 671 79
rect 672 75 676 79
rect 541 49 545 53
rect 546 49 550 53
rect 551 49 555 53
rect 556 49 560 53
rect 541 39 545 43
rect 546 39 550 43
rect 551 39 555 43
rect 556 39 560 43
rect 541 29 545 33
rect 546 29 550 33
rect 551 29 555 33
rect 556 29 560 33
rect 570 49 574 53
rect 575 49 579 53
rect 580 49 584 53
rect 585 49 589 53
rect 570 39 574 43
rect 575 39 579 43
rect 580 39 584 43
rect 585 39 589 43
rect 570 29 574 33
rect 575 29 579 33
rect 580 29 584 33
rect 585 29 589 33
rect 599 49 603 53
rect 604 49 608 53
rect 609 49 613 53
rect 614 49 618 53
rect 599 39 603 43
rect 604 39 608 43
rect 609 39 613 43
rect 614 39 618 43
rect 599 29 603 33
rect 604 29 608 33
rect 609 29 613 33
rect 614 29 618 33
rect 628 49 632 53
rect 633 49 637 53
rect 638 49 642 53
rect 643 49 647 53
rect 628 39 632 43
rect 633 39 637 43
rect 638 39 642 43
rect 643 39 647 43
rect 628 29 632 33
rect 633 29 637 33
rect 638 29 642 33
rect 643 29 647 33
rect 657 49 661 53
rect 662 49 666 53
rect 667 49 671 53
rect 672 49 676 53
rect 657 39 661 43
rect 662 39 666 43
rect 667 39 671 43
rect 672 39 676 43
rect 657 29 661 33
rect 662 29 666 33
rect 667 29 671 33
rect 672 29 676 33
rect 357 -44 361 -40
rect 367 -44 371 -40
rect 377 -44 381 -40
rect 357 -49 361 -45
rect 367 -49 371 -45
rect 377 -49 381 -45
rect 357 -54 361 -50
rect 367 -54 371 -50
rect 377 -54 381 -50
rect 357 -59 361 -55
rect 367 -59 371 -55
rect 377 -59 381 -55
rect 403 -44 407 -40
rect 413 -44 417 -40
rect 423 -44 427 -40
rect 403 -49 407 -45
rect 413 -49 417 -45
rect 423 -49 427 -45
rect 403 -54 407 -50
rect 413 -54 417 -50
rect 423 -54 427 -50
rect 403 -59 407 -55
rect 413 -59 417 -55
rect 423 -59 427 -55
rect 357 -70 361 -66
rect 367 -70 371 -66
rect 377 -70 381 -66
rect 357 -75 361 -71
rect 367 -75 371 -71
rect 377 -75 381 -71
rect 357 -80 361 -76
rect 367 -80 371 -76
rect 377 -80 381 -76
rect 357 -85 361 -81
rect 367 -85 371 -81
rect 377 -85 381 -81
rect 403 -70 407 -66
rect 413 -70 417 -66
rect 423 -70 427 -66
rect 403 -75 407 -71
rect 413 -75 417 -71
rect 423 -75 427 -71
rect 403 -80 407 -76
rect 413 -80 417 -76
rect 423 -80 427 -76
rect 403 -85 407 -81
rect 413 -85 417 -81
rect 423 -85 427 -81
rect 357 -96 361 -92
rect 367 -96 371 -92
rect 377 -96 381 -92
rect 357 -101 361 -97
rect 367 -101 371 -97
rect 377 -101 381 -97
rect 357 -106 361 -102
rect 367 -106 371 -102
rect 377 -106 381 -102
rect 357 -111 361 -107
rect 367 -111 371 -107
rect 377 -111 381 -107
rect 403 -96 407 -92
rect 413 -96 417 -92
rect 423 -96 427 -92
rect 403 -101 407 -97
rect 413 -101 417 -97
rect 423 -101 427 -97
rect 403 -106 407 -102
rect 413 -106 417 -102
rect 423 -106 427 -102
rect 403 -111 407 -107
rect 413 -111 417 -107
rect 423 -111 427 -107
rect 357 -122 361 -118
rect 367 -122 371 -118
rect 377 -122 381 -118
rect 357 -127 361 -123
rect 367 -127 371 -123
rect 377 -127 381 -123
rect 357 -132 361 -128
rect 367 -132 371 -128
rect 377 -132 381 -128
rect 357 -137 361 -133
rect 367 -137 371 -133
rect 377 -137 381 -133
rect 403 -122 407 -118
rect 413 -122 417 -118
rect 423 -122 427 -118
rect 403 -127 407 -123
rect 413 -127 417 -123
rect 423 -127 427 -123
rect 403 -132 407 -128
rect 413 -132 417 -128
rect 423 -132 427 -128
rect 403 -137 407 -133
rect 413 -137 417 -133
rect 423 -137 427 -133
rect 357 -148 361 -144
rect 367 -148 371 -144
rect 377 -148 381 -144
rect 357 -153 361 -149
rect 367 -153 371 -149
rect 377 -153 381 -149
rect 357 -158 361 -154
rect 367 -158 371 -154
rect 377 -158 381 -154
rect 357 -163 361 -159
rect 367 -163 371 -159
rect 377 -163 381 -159
rect 403 -148 407 -144
rect 413 -148 417 -144
rect 423 -148 427 -144
rect 403 -153 407 -149
rect 413 -153 417 -149
rect 423 -153 427 -149
rect 403 -158 407 -154
rect 413 -158 417 -154
rect 423 -158 427 -154
rect 403 -163 407 -159
rect 413 -163 417 -159
rect 423 -163 427 -159
<< metal2 >>
rect -143 124 763 618
rect -143 -314 332 124
rect 545 100 546 104
rect 550 100 551 104
rect 555 100 556 104
rect 541 99 560 100
rect 545 95 546 99
rect 550 95 551 99
rect 555 95 556 99
rect 541 94 560 95
rect 545 90 546 94
rect 550 90 551 94
rect 555 90 556 94
rect 541 89 560 90
rect 545 85 546 89
rect 550 85 551 89
rect 555 85 556 89
rect 541 84 560 85
rect 545 80 546 84
rect 550 80 551 84
rect 555 80 556 84
rect 541 79 560 80
rect 545 75 546 79
rect 550 75 551 79
rect 555 75 556 79
rect 541 74 560 75
rect 545 70 546 74
rect 550 70 551 74
rect 555 70 556 74
rect 574 100 575 104
rect 579 100 580 104
rect 584 100 585 104
rect 570 99 589 100
rect 574 95 575 99
rect 579 95 580 99
rect 584 95 585 99
rect 570 94 589 95
rect 574 90 575 94
rect 579 90 580 94
rect 584 90 585 94
rect 570 89 589 90
rect 574 85 575 89
rect 579 85 580 89
rect 584 85 585 89
rect 570 84 589 85
rect 574 80 575 84
rect 579 80 580 84
rect 584 80 585 84
rect 570 79 589 80
rect 574 75 575 79
rect 579 75 580 79
rect 584 75 585 79
rect 570 74 589 75
rect 574 70 575 74
rect 579 70 580 74
rect 584 70 585 74
rect 603 100 604 104
rect 608 100 609 104
rect 613 100 614 104
rect 599 99 618 100
rect 603 95 604 99
rect 608 95 609 99
rect 613 95 614 99
rect 599 94 618 95
rect 603 90 604 94
rect 608 90 609 94
rect 613 90 614 94
rect 599 89 618 90
rect 603 85 604 89
rect 608 85 609 89
rect 613 85 614 89
rect 599 84 618 85
rect 603 80 604 84
rect 608 80 609 84
rect 613 80 614 84
rect 599 79 618 80
rect 603 75 604 79
rect 608 75 609 79
rect 613 75 614 79
rect 599 74 618 75
rect 603 70 604 74
rect 608 70 609 74
rect 613 70 614 74
rect 632 100 633 104
rect 637 100 638 104
rect 642 100 643 104
rect 628 99 647 100
rect 632 95 633 99
rect 637 95 638 99
rect 642 95 643 99
rect 628 94 647 95
rect 632 90 633 94
rect 637 90 638 94
rect 642 90 643 94
rect 628 89 647 90
rect 632 85 633 89
rect 637 85 638 89
rect 642 85 643 89
rect 628 84 647 85
rect 632 80 633 84
rect 637 80 638 84
rect 642 80 643 84
rect 628 79 647 80
rect 632 75 633 79
rect 637 75 638 79
rect 642 75 643 79
rect 628 74 647 75
rect 632 70 633 74
rect 637 70 638 74
rect 642 70 643 74
rect 661 100 662 104
rect 666 100 667 104
rect 671 100 672 104
rect 657 99 676 100
rect 661 95 662 99
rect 666 95 667 99
rect 671 95 672 99
rect 657 94 676 95
rect 661 90 662 94
rect 666 90 667 94
rect 671 90 672 94
rect 657 89 676 90
rect 661 85 662 89
rect 666 85 667 89
rect 671 85 672 89
rect 657 84 676 85
rect 661 80 662 84
rect 666 80 667 84
rect 671 80 672 84
rect 657 79 676 80
rect 661 75 662 79
rect 666 75 667 79
rect 671 75 672 79
rect 657 74 676 75
rect 661 70 662 74
rect 666 70 667 74
rect 671 70 672 74
rect 545 54 546 58
rect 550 54 551 58
rect 555 54 556 58
rect 541 53 560 54
rect 545 49 546 53
rect 550 49 551 53
rect 555 49 556 53
rect 541 48 560 49
rect 545 44 546 48
rect 550 44 551 48
rect 555 44 556 48
rect 541 43 560 44
rect 545 39 546 43
rect 550 39 551 43
rect 555 39 556 43
rect 541 38 560 39
rect 545 34 546 38
rect 550 34 551 38
rect 555 34 556 38
rect 541 33 560 34
rect 545 29 546 33
rect 550 29 551 33
rect 555 29 556 33
rect 541 28 560 29
rect 545 24 546 28
rect 550 24 551 28
rect 555 24 556 28
rect 574 54 575 58
rect 579 54 580 58
rect 584 54 585 58
rect 570 53 589 54
rect 574 49 575 53
rect 579 49 580 53
rect 584 49 585 53
rect 570 48 589 49
rect 574 44 575 48
rect 579 44 580 48
rect 584 44 585 48
rect 570 43 589 44
rect 574 39 575 43
rect 579 39 580 43
rect 584 39 585 43
rect 570 38 589 39
rect 574 34 575 38
rect 579 34 580 38
rect 584 34 585 38
rect 570 33 589 34
rect 574 29 575 33
rect 579 29 580 33
rect 584 29 585 33
rect 570 28 589 29
rect 574 24 575 28
rect 579 24 580 28
rect 584 24 585 28
rect 603 54 604 58
rect 608 54 609 58
rect 613 54 614 58
rect 599 53 618 54
rect 603 49 604 53
rect 608 49 609 53
rect 613 49 614 53
rect 599 48 618 49
rect 603 44 604 48
rect 608 44 609 48
rect 613 44 614 48
rect 599 43 618 44
rect 603 39 604 43
rect 608 39 609 43
rect 613 39 614 43
rect 599 38 618 39
rect 603 34 604 38
rect 608 34 609 38
rect 613 34 614 38
rect 599 33 618 34
rect 603 29 604 33
rect 608 29 609 33
rect 613 29 614 33
rect 599 28 618 29
rect 603 24 604 28
rect 608 24 609 28
rect 613 24 614 28
rect 632 54 633 58
rect 637 54 638 58
rect 642 54 643 58
rect 628 53 647 54
rect 632 49 633 53
rect 637 49 638 53
rect 642 49 643 53
rect 628 48 647 49
rect 632 44 633 48
rect 637 44 638 48
rect 642 44 643 48
rect 628 43 647 44
rect 632 39 633 43
rect 637 39 638 43
rect 642 39 643 43
rect 628 38 647 39
rect 632 34 633 38
rect 637 34 638 38
rect 642 34 643 38
rect 628 33 647 34
rect 632 29 633 33
rect 637 29 638 33
rect 642 29 643 33
rect 628 28 647 29
rect 632 24 633 28
rect 637 24 638 28
rect 642 24 643 28
rect 661 54 662 58
rect 666 54 667 58
rect 671 54 672 58
rect 657 53 676 54
rect 661 49 662 53
rect 666 49 667 53
rect 671 49 672 53
rect 657 48 676 49
rect 661 44 662 48
rect 666 44 667 48
rect 671 44 672 48
rect 657 43 676 44
rect 661 39 662 43
rect 666 39 667 43
rect 671 39 672 43
rect 657 38 676 39
rect 661 34 662 38
rect 666 34 667 38
rect 671 34 672 38
rect 657 33 676 34
rect 661 29 662 33
rect 666 29 667 33
rect 671 29 672 33
rect 657 28 676 29
rect 661 24 662 28
rect 666 24 667 28
rect 671 24 672 28
rect 356 -44 357 -40
rect 361 -44 362 -40
rect 366 -44 367 -40
rect 371 -44 372 -40
rect 376 -44 377 -40
rect 381 -44 382 -40
rect 352 -45 386 -44
rect 356 -49 357 -45
rect 361 -49 362 -45
rect 366 -49 367 -45
rect 371 -49 372 -45
rect 376 -49 377 -45
rect 381 -49 382 -45
rect 352 -50 386 -49
rect 356 -54 357 -50
rect 361 -54 362 -50
rect 366 -54 367 -50
rect 371 -54 372 -50
rect 376 -54 377 -50
rect 381 -54 382 -50
rect 352 -55 386 -54
rect 356 -59 357 -55
rect 361 -59 362 -55
rect 366 -59 367 -55
rect 371 -59 372 -55
rect 376 -59 377 -55
rect 381 -59 382 -55
rect 402 -44 403 -40
rect 407 -44 408 -40
rect 412 -44 413 -40
rect 417 -44 418 -40
rect 422 -44 423 -40
rect 427 -44 428 -40
rect 398 -45 432 -44
rect 402 -49 403 -45
rect 407 -49 408 -45
rect 412 -49 413 -45
rect 417 -49 418 -45
rect 422 -49 423 -45
rect 427 -49 428 -45
rect 398 -50 432 -49
rect 402 -54 403 -50
rect 407 -54 408 -50
rect 412 -54 413 -50
rect 417 -54 418 -50
rect 422 -54 423 -50
rect 427 -54 428 -50
rect 398 -55 432 -54
rect 402 -59 403 -55
rect 407 -59 408 -55
rect 412 -59 413 -55
rect 417 -59 418 -55
rect 422 -59 423 -55
rect 427 -59 428 -55
rect 356 -70 357 -66
rect 361 -70 362 -66
rect 366 -70 367 -66
rect 371 -70 372 -66
rect 376 -70 377 -66
rect 381 -70 382 -66
rect 352 -71 386 -70
rect 356 -75 357 -71
rect 361 -75 362 -71
rect 366 -75 367 -71
rect 371 -75 372 -71
rect 376 -75 377 -71
rect 381 -75 382 -71
rect 352 -76 386 -75
rect 356 -80 357 -76
rect 361 -80 362 -76
rect 366 -80 367 -76
rect 371 -80 372 -76
rect 376 -80 377 -76
rect 381 -80 382 -76
rect 352 -81 386 -80
rect 356 -85 357 -81
rect 361 -85 362 -81
rect 366 -85 367 -81
rect 371 -85 372 -81
rect 376 -85 377 -81
rect 381 -85 382 -81
rect 402 -70 403 -66
rect 407 -70 408 -66
rect 412 -70 413 -66
rect 417 -70 418 -66
rect 422 -70 423 -66
rect 427 -70 428 -66
rect 398 -71 432 -70
rect 402 -75 403 -71
rect 407 -75 408 -71
rect 412 -75 413 -71
rect 417 -75 418 -71
rect 422 -75 423 -71
rect 427 -75 428 -71
rect 398 -76 432 -75
rect 402 -80 403 -76
rect 407 -80 408 -76
rect 412 -80 413 -76
rect 417 -80 418 -76
rect 422 -80 423 -76
rect 427 -80 428 -76
rect 398 -81 432 -80
rect 402 -85 403 -81
rect 407 -85 408 -81
rect 412 -85 413 -81
rect 417 -85 418 -81
rect 422 -85 423 -81
rect 427 -85 428 -81
rect 356 -96 357 -92
rect 361 -96 362 -92
rect 366 -96 367 -92
rect 371 -96 372 -92
rect 376 -96 377 -92
rect 381 -96 382 -92
rect 352 -97 386 -96
rect 356 -101 357 -97
rect 361 -101 362 -97
rect 366 -101 367 -97
rect 371 -101 372 -97
rect 376 -101 377 -97
rect 381 -101 382 -97
rect 352 -102 386 -101
rect 356 -106 357 -102
rect 361 -106 362 -102
rect 366 -106 367 -102
rect 371 -106 372 -102
rect 376 -106 377 -102
rect 381 -106 382 -102
rect 352 -107 386 -106
rect 356 -111 357 -107
rect 361 -111 362 -107
rect 366 -111 367 -107
rect 371 -111 372 -107
rect 376 -111 377 -107
rect 381 -111 382 -107
rect 402 -96 403 -92
rect 407 -96 408 -92
rect 412 -96 413 -92
rect 417 -96 418 -92
rect 422 -96 423 -92
rect 427 -96 428 -92
rect 398 -97 432 -96
rect 402 -101 403 -97
rect 407 -101 408 -97
rect 412 -101 413 -97
rect 417 -101 418 -97
rect 422 -101 423 -97
rect 427 -101 428 -97
rect 398 -102 432 -101
rect 402 -106 403 -102
rect 407 -106 408 -102
rect 412 -106 413 -102
rect 417 -106 418 -102
rect 422 -106 423 -102
rect 427 -106 428 -102
rect 398 -107 432 -106
rect 402 -111 403 -107
rect 407 -111 408 -107
rect 412 -111 413 -107
rect 417 -111 418 -107
rect 422 -111 423 -107
rect 427 -111 428 -107
rect 356 -122 357 -118
rect 361 -122 362 -118
rect 366 -122 367 -118
rect 371 -122 372 -118
rect 376 -122 377 -118
rect 381 -122 382 -118
rect 352 -123 386 -122
rect 356 -127 357 -123
rect 361 -127 362 -123
rect 366 -127 367 -123
rect 371 -127 372 -123
rect 376 -127 377 -123
rect 381 -127 382 -123
rect 352 -128 386 -127
rect 356 -132 357 -128
rect 361 -132 362 -128
rect 366 -132 367 -128
rect 371 -132 372 -128
rect 376 -132 377 -128
rect 381 -132 382 -128
rect 352 -133 386 -132
rect 356 -137 357 -133
rect 361 -137 362 -133
rect 366 -137 367 -133
rect 371 -137 372 -133
rect 376 -137 377 -133
rect 381 -137 382 -133
rect 402 -122 403 -118
rect 407 -122 408 -118
rect 412 -122 413 -118
rect 417 -122 418 -118
rect 422 -122 423 -118
rect 427 -122 428 -118
rect 398 -123 432 -122
rect 402 -127 403 -123
rect 407 -127 408 -123
rect 412 -127 413 -123
rect 417 -127 418 -123
rect 422 -127 423 -123
rect 427 -127 428 -123
rect 398 -128 432 -127
rect 402 -132 403 -128
rect 407 -132 408 -128
rect 412 -132 413 -128
rect 417 -132 418 -128
rect 422 -132 423 -128
rect 427 -132 428 -128
rect 398 -133 432 -132
rect 402 -137 403 -133
rect 407 -137 408 -133
rect 412 -137 413 -133
rect 417 -137 418 -133
rect 422 -137 423 -133
rect 427 -137 428 -133
rect 356 -148 357 -144
rect 361 -148 362 -144
rect 366 -148 367 -144
rect 371 -148 372 -144
rect 376 -148 377 -144
rect 381 -148 382 -144
rect 352 -149 386 -148
rect 356 -153 357 -149
rect 361 -153 362 -149
rect 366 -153 367 -149
rect 371 -153 372 -149
rect 376 -153 377 -149
rect 381 -153 382 -149
rect 352 -154 386 -153
rect 356 -158 357 -154
rect 361 -158 362 -154
rect 366 -158 367 -154
rect 371 -158 372 -154
rect 376 -158 377 -154
rect 381 -158 382 -154
rect 352 -159 386 -158
rect 356 -163 357 -159
rect 361 -163 362 -159
rect 366 -163 367 -159
rect 371 -163 372 -159
rect 376 -163 377 -159
rect 381 -163 382 -159
rect 402 -148 403 -144
rect 407 -148 408 -144
rect 412 -148 413 -144
rect 417 -148 418 -144
rect 422 -148 423 -144
rect 427 -148 428 -144
rect 398 -149 432 -148
rect 402 -153 403 -149
rect 407 -153 408 -149
rect 412 -153 413 -149
rect 417 -153 418 -149
rect 422 -153 423 -149
rect 427 -153 428 -149
rect 398 -154 432 -153
rect 402 -158 403 -154
rect 407 -158 408 -154
rect 412 -158 413 -154
rect 417 -158 418 -154
rect 422 -158 423 -154
rect 427 -158 428 -154
rect 398 -159 432 -158
rect 402 -163 403 -159
rect 407 -163 408 -159
rect 412 -163 413 -159
rect 417 -163 418 -159
rect 422 -163 423 -159
rect 427 -163 428 -159
<< m3contact >>
rect 541 100 545 104
rect 546 100 550 104
rect 551 100 555 104
rect 556 100 560 104
rect 541 90 545 94
rect 546 90 550 94
rect 551 90 555 94
rect 556 90 560 94
rect 541 80 545 84
rect 546 80 550 84
rect 551 80 555 84
rect 556 80 560 84
rect 541 70 545 74
rect 546 70 550 74
rect 551 70 555 74
rect 556 70 560 74
rect 570 100 574 104
rect 575 100 579 104
rect 580 100 584 104
rect 585 100 589 104
rect 570 90 574 94
rect 575 90 579 94
rect 580 90 584 94
rect 585 90 589 94
rect 570 80 574 84
rect 575 80 579 84
rect 580 80 584 84
rect 585 80 589 84
rect 570 70 574 74
rect 575 70 579 74
rect 580 70 584 74
rect 585 70 589 74
rect 599 100 603 104
rect 604 100 608 104
rect 609 100 613 104
rect 614 100 618 104
rect 599 90 603 94
rect 604 90 608 94
rect 609 90 613 94
rect 614 90 618 94
rect 599 80 603 84
rect 604 80 608 84
rect 609 80 613 84
rect 614 80 618 84
rect 599 70 603 74
rect 604 70 608 74
rect 609 70 613 74
rect 614 70 618 74
rect 628 100 632 104
rect 633 100 637 104
rect 638 100 642 104
rect 643 100 647 104
rect 628 90 632 94
rect 633 90 637 94
rect 638 90 642 94
rect 643 90 647 94
rect 628 80 632 84
rect 633 80 637 84
rect 638 80 642 84
rect 643 80 647 84
rect 628 70 632 74
rect 633 70 637 74
rect 638 70 642 74
rect 643 70 647 74
rect 657 100 661 104
rect 662 100 666 104
rect 667 100 671 104
rect 672 100 676 104
rect 657 90 661 94
rect 662 90 666 94
rect 667 90 671 94
rect 672 90 676 94
rect 657 80 661 84
rect 662 80 666 84
rect 667 80 671 84
rect 672 80 676 84
rect 657 70 661 74
rect 662 70 666 74
rect 667 70 671 74
rect 672 70 676 74
rect 541 54 545 58
rect 546 54 550 58
rect 551 54 555 58
rect 556 54 560 58
rect 541 44 545 48
rect 546 44 550 48
rect 551 44 555 48
rect 556 44 560 48
rect 541 34 545 38
rect 546 34 550 38
rect 551 34 555 38
rect 556 34 560 38
rect 541 24 545 28
rect 546 24 550 28
rect 551 24 555 28
rect 556 24 560 28
rect 570 54 574 58
rect 575 54 579 58
rect 580 54 584 58
rect 585 54 589 58
rect 570 44 574 48
rect 575 44 579 48
rect 580 44 584 48
rect 585 44 589 48
rect 570 34 574 38
rect 575 34 579 38
rect 580 34 584 38
rect 585 34 589 38
rect 570 24 574 28
rect 575 24 579 28
rect 580 24 584 28
rect 585 24 589 28
rect 599 54 603 58
rect 604 54 608 58
rect 609 54 613 58
rect 614 54 618 58
rect 599 44 603 48
rect 604 44 608 48
rect 609 44 613 48
rect 614 44 618 48
rect 599 34 603 38
rect 604 34 608 38
rect 609 34 613 38
rect 614 34 618 38
rect 599 24 603 28
rect 604 24 608 28
rect 609 24 613 28
rect 614 24 618 28
rect 628 54 632 58
rect 633 54 637 58
rect 638 54 642 58
rect 643 54 647 58
rect 628 44 632 48
rect 633 44 637 48
rect 638 44 642 48
rect 643 44 647 48
rect 628 34 632 38
rect 633 34 637 38
rect 638 34 642 38
rect 643 34 647 38
rect 628 24 632 28
rect 633 24 637 28
rect 638 24 642 28
rect 643 24 647 28
rect 657 54 661 58
rect 662 54 666 58
rect 667 54 671 58
rect 672 54 676 58
rect 657 44 661 48
rect 662 44 666 48
rect 667 44 671 48
rect 672 44 676 48
rect 657 34 661 38
rect 662 34 666 38
rect 667 34 671 38
rect 672 34 676 38
rect 657 24 661 28
rect 662 24 666 28
rect 667 24 671 28
rect 672 24 676 28
rect 352 -44 356 -40
rect 362 -44 366 -40
rect 372 -44 376 -40
rect 382 -44 386 -40
rect 352 -49 356 -45
rect 362 -49 366 -45
rect 372 -49 376 -45
rect 382 -49 386 -45
rect 352 -54 356 -50
rect 362 -54 366 -50
rect 372 -54 376 -50
rect 382 -54 386 -50
rect 352 -59 356 -55
rect 362 -59 366 -55
rect 372 -59 376 -55
rect 382 -59 386 -55
rect 398 -44 402 -40
rect 408 -44 412 -40
rect 418 -44 422 -40
rect 428 -44 432 -40
rect 398 -49 402 -45
rect 408 -49 412 -45
rect 418 -49 422 -45
rect 428 -49 432 -45
rect 398 -54 402 -50
rect 408 -54 412 -50
rect 418 -54 422 -50
rect 428 -54 432 -50
rect 398 -59 402 -55
rect 408 -59 412 -55
rect 418 -59 422 -55
rect 428 -59 432 -55
rect 352 -70 356 -66
rect 362 -70 366 -66
rect 372 -70 376 -66
rect 382 -70 386 -66
rect 352 -75 356 -71
rect 362 -75 366 -71
rect 372 -75 376 -71
rect 382 -75 386 -71
rect 352 -80 356 -76
rect 362 -80 366 -76
rect 372 -80 376 -76
rect 382 -80 386 -76
rect 352 -85 356 -81
rect 362 -85 366 -81
rect 372 -85 376 -81
rect 382 -85 386 -81
rect 398 -70 402 -66
rect 408 -70 412 -66
rect 418 -70 422 -66
rect 428 -70 432 -66
rect 398 -75 402 -71
rect 408 -75 412 -71
rect 418 -75 422 -71
rect 428 -75 432 -71
rect 398 -80 402 -76
rect 408 -80 412 -76
rect 418 -80 422 -76
rect 428 -80 432 -76
rect 398 -85 402 -81
rect 408 -85 412 -81
rect 418 -85 422 -81
rect 428 -85 432 -81
rect 352 -96 356 -92
rect 362 -96 366 -92
rect 372 -96 376 -92
rect 382 -96 386 -92
rect 352 -101 356 -97
rect 362 -101 366 -97
rect 372 -101 376 -97
rect 382 -101 386 -97
rect 352 -106 356 -102
rect 362 -106 366 -102
rect 372 -106 376 -102
rect 382 -106 386 -102
rect 352 -111 356 -107
rect 362 -111 366 -107
rect 372 -111 376 -107
rect 382 -111 386 -107
rect 398 -96 402 -92
rect 408 -96 412 -92
rect 418 -96 422 -92
rect 428 -96 432 -92
rect 398 -101 402 -97
rect 408 -101 412 -97
rect 418 -101 422 -97
rect 428 -101 432 -97
rect 398 -106 402 -102
rect 408 -106 412 -102
rect 418 -106 422 -102
rect 428 -106 432 -102
rect 398 -111 402 -107
rect 408 -111 412 -107
rect 418 -111 422 -107
rect 428 -111 432 -107
rect 352 -122 356 -118
rect 362 -122 366 -118
rect 372 -122 376 -118
rect 382 -122 386 -118
rect 352 -127 356 -123
rect 362 -127 366 -123
rect 372 -127 376 -123
rect 382 -127 386 -123
rect 352 -132 356 -128
rect 362 -132 366 -128
rect 372 -132 376 -128
rect 382 -132 386 -128
rect 352 -137 356 -133
rect 362 -137 366 -133
rect 372 -137 376 -133
rect 382 -137 386 -133
rect 398 -122 402 -118
rect 408 -122 412 -118
rect 418 -122 422 -118
rect 428 -122 432 -118
rect 398 -127 402 -123
rect 408 -127 412 -123
rect 418 -127 422 -123
rect 428 -127 432 -123
rect 398 -132 402 -128
rect 408 -132 412 -128
rect 418 -132 422 -128
rect 428 -132 432 -128
rect 398 -137 402 -133
rect 408 -137 412 -133
rect 418 -137 422 -133
rect 428 -137 432 -133
rect 352 -148 356 -144
rect 362 -148 366 -144
rect 372 -148 376 -144
rect 382 -148 386 -144
rect 352 -153 356 -149
rect 362 -153 366 -149
rect 372 -153 376 -149
rect 382 -153 386 -149
rect 352 -158 356 -154
rect 362 -158 366 -154
rect 372 -158 376 -154
rect 382 -158 386 -154
rect 352 -163 356 -159
rect 362 -163 366 -159
rect 372 -163 376 -159
rect 382 -163 386 -159
rect 398 -148 402 -144
rect 408 -148 412 -144
rect 418 -148 422 -144
rect 428 -148 432 -144
rect 398 -153 402 -149
rect 408 -153 412 -149
rect 418 -153 422 -149
rect 428 -153 432 -149
rect 398 -158 402 -154
rect 408 -158 412 -154
rect 418 -158 422 -154
rect 428 -158 432 -154
rect 398 -163 402 -159
rect 408 -163 412 -159
rect 418 -163 422 -159
rect 428 -163 432 -159
<< metal3 >>
rect 309 104 774 147
rect 309 100 541 104
rect 545 100 546 104
rect 550 100 551 104
rect 555 100 556 104
rect 560 100 570 104
rect 574 100 575 104
rect 579 100 580 104
rect 584 100 585 104
rect 589 100 599 104
rect 603 100 604 104
rect 608 100 609 104
rect 613 100 614 104
rect 618 100 628 104
rect 632 100 633 104
rect 637 100 638 104
rect 642 100 643 104
rect 647 100 657 104
rect 661 100 662 104
rect 666 100 667 104
rect 671 100 672 104
rect 676 100 774 104
rect 309 94 774 100
rect 309 90 541 94
rect 545 90 546 94
rect 550 90 551 94
rect 555 90 556 94
rect 560 90 570 94
rect 574 90 575 94
rect 579 90 580 94
rect 584 90 585 94
rect 589 90 599 94
rect 603 90 604 94
rect 608 90 609 94
rect 613 90 614 94
rect 618 90 628 94
rect 632 90 633 94
rect 637 90 638 94
rect 642 90 643 94
rect 647 90 657 94
rect 661 90 662 94
rect 666 90 667 94
rect 671 90 672 94
rect 676 90 774 94
rect 309 84 774 90
rect 309 80 541 84
rect 545 80 546 84
rect 550 80 551 84
rect 555 80 556 84
rect 560 80 570 84
rect 574 80 575 84
rect 579 80 580 84
rect 584 80 585 84
rect 589 80 599 84
rect 603 80 604 84
rect 608 80 609 84
rect 613 80 614 84
rect 618 80 628 84
rect 632 80 633 84
rect 637 80 638 84
rect 642 80 643 84
rect 647 80 657 84
rect 661 80 662 84
rect 666 80 667 84
rect 671 80 672 84
rect 676 80 774 84
rect 309 74 774 80
rect 309 70 541 74
rect 545 70 546 74
rect 550 70 551 74
rect 555 70 556 74
rect 560 70 570 74
rect 574 70 575 74
rect 579 70 580 74
rect 584 70 585 74
rect 589 70 599 74
rect 603 70 604 74
rect 608 70 609 74
rect 613 70 614 74
rect 618 70 628 74
rect 632 70 633 74
rect 637 70 638 74
rect 642 70 643 74
rect 647 70 657 74
rect 661 70 662 74
rect 666 70 667 74
rect 671 70 672 74
rect 676 70 774 74
rect 309 67 774 70
rect 309 -40 389 67
rect 309 -44 352 -40
rect 356 -44 362 -40
rect 366 -44 372 -40
rect 376 -44 382 -40
rect 386 -44 389 -40
rect 309 -45 389 -44
rect 309 -49 352 -45
rect 356 -49 362 -45
rect 366 -49 372 -45
rect 376 -49 382 -45
rect 386 -49 389 -45
rect 309 -50 389 -49
rect 309 -54 352 -50
rect 356 -54 362 -50
rect 366 -54 372 -50
rect 376 -54 382 -50
rect 386 -54 389 -50
rect 309 -55 389 -54
rect 309 -59 352 -55
rect 356 -59 362 -55
rect 366 -59 372 -55
rect 376 -59 382 -55
rect 386 -59 389 -55
rect 309 -66 389 -59
rect 309 -70 352 -66
rect 356 -70 362 -66
rect 366 -70 372 -66
rect 376 -70 382 -66
rect 386 -70 389 -66
rect 309 -71 389 -70
rect 309 -75 352 -71
rect 356 -75 362 -71
rect 366 -75 372 -71
rect 376 -75 382 -71
rect 386 -75 389 -71
rect 309 -76 389 -75
rect 309 -80 352 -76
rect 356 -80 362 -76
rect 366 -80 372 -76
rect 376 -80 382 -76
rect 386 -80 389 -76
rect 309 -81 389 -80
rect 309 -85 352 -81
rect 356 -85 362 -81
rect 366 -85 372 -81
rect 376 -85 382 -81
rect 386 -85 389 -81
rect 309 -92 389 -85
rect 309 -96 352 -92
rect 356 -96 362 -92
rect 366 -96 372 -92
rect 376 -96 382 -92
rect 386 -96 389 -92
rect 309 -97 389 -96
rect 309 -101 352 -97
rect 356 -101 362 -97
rect 366 -101 372 -97
rect 376 -101 382 -97
rect 386 -101 389 -97
rect 309 -102 389 -101
rect 309 -106 352 -102
rect 356 -106 362 -102
rect 366 -106 372 -102
rect 376 -106 382 -102
rect 386 -106 389 -102
rect 309 -107 389 -106
rect 309 -111 352 -107
rect 356 -111 362 -107
rect 366 -111 372 -107
rect 376 -111 382 -107
rect 386 -111 389 -107
rect 309 -118 389 -111
rect 309 -122 352 -118
rect 356 -122 362 -118
rect 366 -122 372 -118
rect 376 -122 382 -118
rect 386 -122 389 -118
rect 309 -123 389 -122
rect 309 -127 352 -123
rect 356 -127 362 -123
rect 366 -127 372 -123
rect 376 -127 382 -123
rect 386 -127 389 -123
rect 309 -128 389 -127
rect 309 -132 352 -128
rect 356 -132 362 -128
rect 366 -132 372 -128
rect 376 -132 382 -128
rect 386 -132 389 -128
rect 309 -133 389 -132
rect 309 -137 352 -133
rect 356 -137 362 -133
rect 366 -137 372 -133
rect 376 -137 382 -133
rect 386 -137 389 -133
rect 309 -144 389 -137
rect 309 -148 352 -144
rect 356 -148 362 -144
rect 366 -148 372 -144
rect 376 -148 382 -144
rect 386 -148 389 -144
rect 309 -149 389 -148
rect 309 -153 352 -149
rect 356 -153 362 -149
rect 366 -153 372 -149
rect 376 -153 382 -149
rect 386 -153 389 -149
rect 309 -154 389 -153
rect 309 -158 352 -154
rect 356 -158 362 -154
rect 366 -158 372 -154
rect 376 -158 382 -154
rect 386 -158 389 -154
rect 309 -159 389 -158
rect 309 -163 352 -159
rect 356 -163 362 -159
rect 366 -163 372 -159
rect 376 -163 382 -159
rect 386 -163 389 -159
rect 309 -331 389 -163
rect 393 58 774 63
rect 393 54 541 58
rect 545 54 546 58
rect 550 54 551 58
rect 555 54 556 58
rect 560 54 570 58
rect 574 54 575 58
rect 579 54 580 58
rect 584 54 585 58
rect 589 54 599 58
rect 603 54 604 58
rect 608 54 609 58
rect 613 54 614 58
rect 618 54 628 58
rect 632 54 633 58
rect 637 54 638 58
rect 642 54 643 58
rect 647 54 657 58
rect 661 54 662 58
rect 666 54 667 58
rect 671 54 672 58
rect 676 54 774 58
rect 393 48 774 54
rect 393 44 541 48
rect 545 44 546 48
rect 550 44 551 48
rect 555 44 556 48
rect 560 44 570 48
rect 574 44 575 48
rect 579 44 580 48
rect 584 44 585 48
rect 589 44 599 48
rect 603 44 604 48
rect 608 44 609 48
rect 613 44 614 48
rect 618 44 628 48
rect 632 44 633 48
rect 637 44 638 48
rect 642 44 643 48
rect 647 44 657 48
rect 661 44 662 48
rect 666 44 667 48
rect 671 44 672 48
rect 676 44 774 48
rect 393 38 774 44
rect 393 34 541 38
rect 545 34 546 38
rect 550 34 551 38
rect 555 34 556 38
rect 560 34 570 38
rect 574 34 575 38
rect 579 34 580 38
rect 584 34 585 38
rect 589 34 599 38
rect 603 34 604 38
rect 608 34 609 38
rect 613 34 614 38
rect 618 34 628 38
rect 632 34 633 38
rect 637 34 638 38
rect 642 34 643 38
rect 647 34 657 38
rect 661 34 662 38
rect 666 34 667 38
rect 671 34 672 38
rect 676 34 774 38
rect 393 28 774 34
rect 393 24 541 28
rect 545 24 546 28
rect 550 24 551 28
rect 555 24 556 28
rect 560 24 570 28
rect 574 24 575 28
rect 579 24 580 28
rect 584 24 585 28
rect 589 24 599 28
rect 603 24 604 28
rect 608 24 609 28
rect 613 24 614 28
rect 618 24 628 28
rect 632 24 633 28
rect 637 24 638 28
rect 642 24 643 28
rect 647 24 657 28
rect 661 24 662 28
rect 666 24 667 28
rect 671 24 672 28
rect 676 24 774 28
rect 393 -40 774 24
rect 393 -44 398 -40
rect 402 -44 408 -40
rect 412 -44 418 -40
rect 422 -44 428 -40
rect 432 -44 774 -40
rect 393 -45 774 -44
rect 393 -49 398 -45
rect 402 -49 408 -45
rect 412 -49 418 -45
rect 422 -49 428 -45
rect 432 -49 774 -45
rect 393 -50 774 -49
rect 393 -54 398 -50
rect 402 -54 408 -50
rect 412 -54 418 -50
rect 422 -54 428 -50
rect 432 -52 774 -50
rect 432 -54 508 -52
rect 393 -55 508 -54
rect 393 -59 398 -55
rect 402 -59 408 -55
rect 412 -59 418 -55
rect 422 -59 428 -55
rect 432 -59 508 -55
rect 393 -66 508 -59
rect 393 -70 398 -66
rect 402 -70 408 -66
rect 412 -70 418 -66
rect 422 -70 428 -66
rect 432 -70 508 -66
rect 393 -71 508 -70
rect 393 -75 398 -71
rect 402 -75 408 -71
rect 412 -75 418 -71
rect 422 -75 428 -71
rect 432 -75 508 -71
rect 393 -76 508 -75
rect 393 -80 398 -76
rect 402 -80 408 -76
rect 412 -80 418 -76
rect 422 -80 428 -76
rect 432 -80 508 -76
rect 393 -81 508 -80
rect 393 -85 398 -81
rect 402 -85 408 -81
rect 412 -85 418 -81
rect 422 -85 428 -81
rect 432 -85 508 -81
rect 393 -92 508 -85
rect 393 -96 398 -92
rect 402 -96 408 -92
rect 412 -96 418 -92
rect 422 -96 428 -92
rect 432 -96 508 -92
rect 393 -97 508 -96
rect 393 -101 398 -97
rect 402 -101 408 -97
rect 412 -101 418 -97
rect 422 -101 428 -97
rect 432 -101 508 -97
rect 393 -102 508 -101
rect 393 -106 398 -102
rect 402 -106 408 -102
rect 412 -106 418 -102
rect 422 -106 428 -102
rect 432 -106 508 -102
rect 393 -107 508 -106
rect 393 -111 398 -107
rect 402 -111 408 -107
rect 412 -111 418 -107
rect 422 -111 428 -107
rect 432 -111 508 -107
rect 393 -118 508 -111
rect 393 -122 398 -118
rect 402 -122 408 -118
rect 412 -122 418 -118
rect 422 -122 428 -118
rect 432 -122 508 -118
rect 393 -123 508 -122
rect 393 -127 398 -123
rect 402 -127 408 -123
rect 412 -127 418 -123
rect 422 -127 428 -123
rect 432 -127 508 -123
rect 393 -128 508 -127
rect 393 -132 398 -128
rect 402 -132 408 -128
rect 412 -132 418 -128
rect 422 -132 428 -128
rect 432 -132 508 -128
rect 393 -133 508 -132
rect 393 -137 398 -133
rect 402 -137 408 -133
rect 412 -137 418 -133
rect 422 -137 428 -133
rect 432 -137 508 -133
rect 393 -144 508 -137
rect 393 -148 398 -144
rect 402 -148 408 -144
rect 412 -148 418 -144
rect 422 -148 428 -144
rect 432 -148 508 -144
rect 393 -149 508 -148
rect 393 -153 398 -149
rect 402 -153 408 -149
rect 412 -153 418 -149
rect 422 -153 428 -149
rect 432 -153 508 -149
rect 393 -154 508 -153
rect 393 -158 398 -154
rect 402 -158 408 -154
rect 412 -158 418 -154
rect 422 -158 428 -154
rect 432 -158 508 -154
rect 393 -159 508 -158
rect 393 -163 398 -159
rect 402 -163 408 -159
rect 412 -163 418 -159
rect 422 -163 428 -159
rect 432 -163 508 -159
rect 393 -331 508 -163
rect 458 -333 508 -331
<< labels >>
rlabel metal3 479 78 479 78 1 Vdd!
rlabel metal3 478 52 478 52 1 GND!
rlabel metal3 378 -317 378 -317 7 Vdd!
rlabel metal3 404 -318 404 -318 7 GND!
<< end >>
