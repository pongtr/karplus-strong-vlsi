magic
tech scmos
timestamp 1512627054
<< nwell >>
rect -35 1319 92 1339
<< pwell >>
rect -49 1290 81 1310
<< ntransistor >>
rect -22 1296 -20 1303
rect -4 1296 -2 1303
rect 14 1296 16 1303
rect 32 1296 34 1303
rect 49 1296 51 1303
rect 68 1296 70 1303
<< ptransistor >>
rect -22 1326 -20 1333
rect -4 1326 -2 1333
rect 14 1326 16 1333
rect 32 1326 34 1333
rect 49 1326 51 1333
rect 68 1326 70 1333
<< ndiffusion >>
rect -28 1301 -22 1303
rect -23 1296 -22 1301
rect -20 1298 -19 1303
rect -20 1296 -14 1298
rect -5 1298 -4 1303
rect -10 1296 -4 1298
rect -2 1298 -1 1303
rect -2 1296 4 1298
rect 8 1301 14 1303
rect 13 1296 14 1301
rect 16 1298 17 1303
rect 16 1296 22 1298
rect 26 1301 32 1303
rect 31 1296 32 1301
rect 34 1298 35 1303
rect 40 1298 49 1303
rect 34 1296 49 1298
rect 51 1298 54 1303
rect 51 1296 59 1298
rect 67 1299 68 1303
rect 63 1296 68 1299
rect 70 1299 71 1303
rect 70 1296 75 1299
<< pdiffusion >>
rect -23 1328 -22 1333
rect -28 1326 -22 1328
rect -20 1331 -14 1333
rect -20 1326 -19 1331
rect -10 1331 -4 1333
rect -5 1326 -4 1331
rect -2 1331 4 1333
rect -2 1326 -1 1331
rect 13 1328 14 1333
rect 8 1326 14 1328
rect 16 1331 22 1333
rect 16 1326 17 1331
rect 31 1328 32 1333
rect 26 1326 32 1328
rect 34 1331 49 1333
rect 34 1326 35 1331
rect 40 1326 49 1331
rect 51 1331 59 1333
rect 51 1326 54 1331
rect 63 1330 68 1333
rect 67 1326 68 1330
rect 70 1330 75 1333
rect 70 1326 71 1330
<< ndcontact >>
rect -28 1296 -23 1301
rect -19 1298 -14 1303
rect -10 1298 -5 1303
rect -1 1298 4 1303
rect 8 1296 13 1301
rect 17 1298 22 1303
rect 26 1296 31 1301
rect 35 1298 40 1303
rect 54 1298 59 1303
rect 63 1299 67 1303
rect 71 1299 75 1303
<< pdcontact >>
rect -28 1328 -23 1333
rect -19 1326 -14 1331
rect -10 1326 -5 1331
rect -1 1326 4 1331
rect 8 1328 13 1333
rect 17 1326 22 1331
rect 26 1328 31 1333
rect 35 1326 40 1331
rect 54 1326 59 1331
rect 63 1326 67 1330
rect 71 1326 75 1330
<< psubstratepcontact >>
rect -46 1297 -41 1302
<< nsubstratencontact >>
rect 80 1327 85 1332
<< polysilicon >>
rect -22 1333 -20 1335
rect -4 1333 -2 1335
rect 14 1333 16 1335
rect 32 1333 34 1335
rect 49 1333 51 1335
rect 68 1333 70 1335
rect -22 1303 -20 1326
rect -4 1324 -2 1326
rect -4 1303 -2 1305
rect 14 1303 16 1326
rect 32 1303 34 1326
rect 49 1325 51 1326
rect 68 1324 70 1326
rect 49 1314 51 1321
rect 49 1312 70 1314
rect 49 1303 51 1305
rect 68 1303 70 1312
rect -22 1294 -20 1296
rect -4 1294 -2 1296
rect 14 1294 16 1296
rect 32 1294 34 1296
rect 49 1291 51 1296
rect 68 1294 70 1296
<< polycontact >>
rect -6 1335 -2 1339
rect 66 1335 70 1339
rect -26 1315 -22 1319
rect 10 1313 14 1317
rect 28 1316 32 1320
rect 47 1321 51 1325
rect -6 1290 -2 1294
rect 47 1287 51 1291
<< metal1 >>
rect -46 1351 -43 1373
rect -46 1348 31 1351
rect -46 1302 -43 1348
rect -28 1333 -23 1348
rect -19 1335 -6 1339
rect -19 1331 -14 1335
rect 8 1333 13 1348
rect -35 1319 -31 1321
rect -40 1315 -26 1319
rect -46 1249 -43 1297
rect -35 1294 -31 1315
rect -19 1303 -14 1326
rect -35 1249 -31 1290
rect -28 1275 -23 1296
rect -10 1312 -5 1326
rect -6 1308 -5 1312
rect -10 1303 -5 1308
rect 26 1333 31 1348
rect -1 1317 4 1326
rect 82 1332 85 1373
rect 17 1320 22 1326
rect -1 1313 10 1317
rect -1 1303 4 1313
rect 10 1309 14 1313
rect 17 1316 28 1320
rect 17 1303 22 1316
rect -19 1287 -14 1298
rect 35 1303 40 1326
rect 8 1275 13 1296
rect 54 1309 59 1326
rect 63 1316 67 1326
rect 63 1309 67 1312
rect 58 1305 67 1309
rect 54 1303 59 1305
rect 63 1303 67 1305
rect 71 1316 75 1326
rect 71 1303 75 1312
rect 26 1275 31 1296
rect 82 1275 85 1327
rect -28 1272 85 1275
rect 82 1249 85 1272
<< m2contact >>
rect -35 1369 -31 1373
rect -2 1335 2 1339
rect -35 1321 -31 1325
rect -35 1290 -31 1294
rect -10 1308 -6 1312
rect 62 1335 66 1339
rect 10 1305 14 1309
rect 25 1312 29 1316
rect 43 1321 47 1325
rect -10 1290 -6 1294
rect -19 1283 -14 1287
rect 63 1312 67 1316
rect 54 1305 58 1309
rect 71 1312 75 1316
rect 47 1283 51 1287
<< metal2 >>
rect -35 1325 -31 1369
rect 2 1335 62 1339
rect 66 1335 70 1339
rect -31 1321 43 1325
rect 29 1312 45 1316
rect 49 1312 63 1316
rect 75 1312 87 1316
rect -40 1308 -10 1312
rect 14 1305 54 1309
rect -31 1290 -10 1294
rect -14 1283 47 1287
<< m3contact >>
rect 87 1312 92 1316
<< metal3 >>
rect 86 1316 93 1317
rect 86 1312 87 1316
rect 92 1312 93 1316
rect 86 1311 93 1312
<< labels >>
rlabel metal1 -39 1349 -39 1349 5 Vdd!
rlabel metal2 -39 1310 -39 1310 1 in
rlabel metal1 -39 1317 -39 1317 1 CLK
rlabel metal1 -16 1317 -16 1317 1 CLKn
rlabel metal2 77 1314 77 1314 1 out
rlabel metal1 81 1273 81 1273 8 GND!
<< end >>
