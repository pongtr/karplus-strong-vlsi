magic
tech scmos
timestamp 1512636464
<< metal1 >>
rect 23 15 27 31
rect 31 11 35 33
rect 39 15 43 28
<< m2contact >>
rect 5 6 9 10
<< metal2 >>
rect 9 6 27 10
use and  and_0
timestamp 1512533720
transform 1 0 -65 0 1 37
box 53 -9 111 29
use stat  stat_0
timestamp 1512532515
transform 1 0 6 0 -1 14
box -3 -7 57 28
<< end >>
