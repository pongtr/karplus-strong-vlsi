magic
tech scmos
timestamp 1512383252
<< nwell >>
rect -5 91 12 95
rect -6 73 12 91
rect 0 11 12 47
rect 0 -33 12 -15
<< pwell >>
rect -6 47 12 73
rect -6 -15 12 11
<< psubstratepcontact >>
rect 2 59 6 63
rect 3 -6 7 -2
<< nsubstratencontact >>
rect 3 28 7 32
rect 3 -25 7 -21
<< metal1 >>
rect 3 70 6 92
rect 3 32 6 52
rect 3 5 6 28
rect 0 1 3 5
rect 3 -21 6 -15
rect 3 -29 6 -25
rect 0 -32 6 -29
<< m2contact >>
rect 3 66 7 70
rect -2 59 2 63
rect 3 52 7 56
rect 3 1 7 5
rect -1 -6 3 -2
rect 3 -15 7 -11
<< metal2 >>
rect 7 66 9 70
rect -6 59 -2 63
rect 6 56 9 66
rect 7 52 9 56
rect -6 -6 -1 -2
rect 7 -15 10 5
rect 0 -25 15 -21
<< end >>
