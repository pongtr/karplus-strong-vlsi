magic
tech scmos
timestamp 1512714235
<< pwell >>
rect -1553 -169 -1540 -157
<< polysilicon >>
rect 1020 1467 1022 1468
rect 988 1445 1012 1447
rect 446 1410 448 1411
rect 418 1388 438 1390
rect -1349 1182 -1347 1189
rect -1212 1182 -1210 1190
rect -1052 1182 -1050 1190
rect -836 1182 -834 1190
rect -508 1182 -506 1190
rect -1563 -89 -1561 -88
rect 1649 -99 1651 -98
rect -1553 -110 -1537 -108
rect 1625 -120 1641 -118
<< polycontact >>
rect 1019 1468 1023 1472
rect 984 1444 988 1448
rect 445 1411 449 1415
rect 414 1387 418 1391
rect 1043 1377 1047 1381
rect 1079 1377 1083 1381
rect 106 1252 110 1256
rect 306 1252 310 1256
rect 499 1251 503 1255
rect 535 1251 539 1255
rect 810 1238 814 1242
rect 810 1229 814 1233
rect -1351 1176 -1345 1182
rect -1214 1176 -1208 1182
rect -1054 1176 -1048 1182
rect -838 1176 -832 1182
rect -510 1176 -504 1182
rect 314 1178 318 1182
rect 810 1114 814 1118
rect 810 1105 814 1109
rect 810 990 814 994
rect 810 981 814 985
rect 810 866 814 870
rect 810 857 814 861
rect 810 742 814 746
rect 810 733 814 737
rect 810 618 814 622
rect 810 609 814 613
rect 810 494 814 498
rect 810 485 814 489
rect 810 370 814 374
rect 810 361 814 365
rect 810 246 814 250
rect 810 237 814 241
rect 810 122 814 126
rect 810 113 814 117
rect -1564 -88 -1560 -84
rect 1648 -98 1652 -94
rect -1537 -111 -1533 -107
rect 1621 -121 1625 -117
rect -1559 -228 -1555 -224
rect -1523 -228 -1519 -224
rect 1650 -226 1654 -222
rect 1686 -226 1690 -222
rect -466 -1462 -462 -1458
rect -458 -1461 -454 -1457
rect 1580 -1462 1584 -1458
rect 1588 -1462 1592 -1458
<< metal1 >>
rect -1481 2331 -1356 2426
rect -1155 2333 -1030 2428
rect -813 2330 -741 2406
rect -503 2335 -431 2411
rect -222 2334 -97 2429
rect 395 2340 520 2435
rect 679 2337 804 2432
rect 1013 2337 1138 2432
rect 1314 2349 1439 2444
rect -2425 1325 -2330 1454
rect -1395 1453 -1382 2007
rect -1116 1817 -1059 1834
rect -1817 1380 -1757 1393
rect -2422 1028 -2327 1157
rect -1817 1071 -1764 1084
rect -2411 685 -2316 814
rect -1817 774 -1776 775
rect -1817 762 -1771 774
rect -2395 378 -2300 507
rect -1818 453 -1778 466
rect -2408 80 -2313 209
rect -1817 144 -1785 157
rect -2406 -250 -2311 -121
rect -1817 -165 -1792 -152
rect -2417 -548 -2322 -419
rect -1817 -474 -1799 -461
rect -2418 -860 -2323 -731
rect -1817 -784 -1806 -769
rect -2406 -1146 -2311 -1017
rect -1817 -1279 -1813 -1079
rect -1810 -1155 -1806 -784
rect -1803 -1031 -1799 -474
rect -1796 -907 -1792 -165
rect -1789 -783 -1785 144
rect -1782 -659 -1778 453
rect -1775 -535 -1771 762
rect -1768 -411 -1764 1071
rect -1761 -287 -1757 1380
rect -1118 1355 -1059 1817
rect -782 1441 -769 2007
rect -781 1363 -769 1441
rect -473 1393 -460 1817
rect -770 1358 -769 1363
rect -188 1322 -134 1819
rect 31 1367 39 1504
rect 31 1363 33 1367
rect 37 1363 39 1367
rect 31 1322 39 1363
rect 43 1360 46 1504
rect 51 1398 54 1504
rect 192 1398 195 1499
rect 51 1395 71 1398
rect 175 1395 195 1398
rect 200 1360 203 1499
rect 43 1357 71 1360
rect 175 1357 203 1360
rect 43 1349 46 1357
rect 200 1354 203 1357
rect 207 1391 215 1499
rect 207 1387 209 1391
rect 213 1387 215 1391
rect 207 1336 215 1387
rect 262 1330 266 1470
rect 445 1415 449 1465
rect 454 1447 467 1817
rect 763 1433 776 1817
rect 1072 1644 1085 1818
rect 1381 1817 1393 1819
rect 1381 1758 1394 1817
rect 810 1637 1085 1644
rect 810 1461 817 1637
rect 992 1407 1017 1411
rect 1065 1407 1071 1411
rect 1081 1396 1084 1406
rect 1065 1393 1084 1396
rect 1043 1381 1047 1393
rect 1095 1381 1099 1390
rect 1090 1377 1099 1381
rect 1103 1381 1107 1394
rect 1119 1377 1123 1406
rect 425 1354 429 1375
rect 429 1350 443 1354
rect 491 1350 501 1354
rect 497 1322 501 1350
rect 504 1336 508 1348
rect 511 1322 515 1332
rect -1637 1304 835 1322
rect -1637 186 -1634 1304
rect -1637 -145 -1634 163
rect -1509 -104 -1506 1261
rect -1376 1245 -1373 1304
rect -1280 1254 -1277 1262
rect -1274 1251 -1270 1304
rect -1266 1257 -1262 1275
rect -1311 1246 -1307 1249
rect -1304 1246 -1300 1249
rect -1297 1246 -1293 1249
rect -1290 1246 -1286 1249
rect -1239 1245 -1236 1304
rect -1143 1255 -1140 1262
rect -1136 1252 -1133 1304
rect -1174 1247 -1170 1250
rect -1167 1247 -1163 1250
rect -1160 1247 -1156 1250
rect -1153 1247 -1149 1250
rect -1079 1245 -1076 1304
rect -983 1255 -980 1262
rect -976 1253 -973 1304
rect -927 1255 -924 1262
rect -863 1245 -860 1304
rect -767 1255 -764 1262
rect -760 1253 -757 1304
rect -535 1245 -532 1304
rect -517 1252 -513 1294
rect -439 1255 -436 1262
rect -432 1253 -429 1304
rect -1516 -108 -1506 -104
rect -1516 -145 -1512 -108
rect -1637 -149 -1606 -145
rect -1554 -149 -1512 -145
rect -1351 -140 -1345 1176
rect -1214 -132 -1208 1176
rect -1054 -124 -1048 1176
rect -838 -116 -832 1176
rect -510 -108 -504 1176
rect -497 -95 -491 1163
rect -484 -82 -478 1171
rect -484 -87 -314 -82
rect -497 -100 -327 -95
rect -510 -113 -340 -108
rect -838 -121 -353 -116
rect -1054 -129 -366 -124
rect -1214 -137 -379 -132
rect -1351 -145 -392 -140
rect -1351 -146 -916 -145
rect -1637 -166 -1634 -149
rect -1559 -163 -1532 -160
rect -1637 -224 -1634 -170
rect -1559 -224 -1555 -163
rect -1516 -190 -1512 -149
rect -1520 -194 -1512 -190
rect -1637 -230 -1563 -224
rect -1536 -224 -1532 -198
rect -1516 -222 -1512 -194
rect -1536 -228 -1523 -224
rect -527 -225 -524 -222
rect -1496 -233 -1492 -229
rect -1489 -233 -1485 -229
rect -1482 -233 -1478 -229
rect -1475 -233 -1471 -229
rect -1468 -233 -1464 -229
rect -1461 -233 -1457 -229
rect -1454 -233 -1450 -229
rect -1447 -233 -1443 -229
rect -1440 -233 -1436 -229
rect -1496 -357 -1492 -353
rect -1489 -357 -1485 -353
rect -1482 -357 -1478 -353
rect -1475 -357 -1471 -353
rect -1468 -357 -1464 -353
rect -1461 -357 -1457 -353
rect -1454 -357 -1450 -353
rect -1447 -357 -1443 -353
rect -1433 -357 -1429 -353
rect -1496 -481 -1492 -477
rect -1489 -481 -1485 -477
rect -1482 -481 -1478 -477
rect -1475 -481 -1471 -477
rect -1468 -481 -1464 -477
rect -1461 -481 -1457 -477
rect -1454 -481 -1450 -477
rect -1440 -481 -1436 -477
rect -1433 -481 -1429 -477
rect -1496 -605 -1492 -601
rect -1489 -605 -1485 -601
rect -1482 -605 -1478 -601
rect -1475 -605 -1471 -601
rect -1468 -605 -1464 -601
rect -1461 -605 -1457 -601
rect -1447 -605 -1443 -601
rect -1440 -605 -1436 -601
rect -1433 -605 -1429 -601
rect -1496 -729 -1492 -725
rect -1489 -729 -1485 -725
rect -1482 -729 -1478 -725
rect -1475 -729 -1471 -725
rect -1468 -729 -1464 -725
rect -1454 -729 -1450 -725
rect -1447 -729 -1443 -725
rect -1440 -729 -1436 -725
rect -1433 -729 -1429 -725
rect -1496 -853 -1492 -849
rect -1489 -853 -1485 -849
rect -1482 -853 -1478 -849
rect -1475 -853 -1471 -849
rect -1454 -853 -1450 -849
rect -1447 -853 -1443 -849
rect -1440 -853 -1436 -849
rect -1433 -853 -1429 -849
rect -1496 -977 -1492 -973
rect -1489 -977 -1485 -973
rect -1482 -977 -1478 -973
rect -1461 -977 -1457 -973
rect -1454 -977 -1450 -973
rect -1447 -977 -1443 -973
rect -1440 -977 -1436 -973
rect -1433 -977 -1429 -973
rect -1496 -1101 -1492 -1097
rect -1489 -1101 -1485 -1097
rect -1468 -1101 -1464 -1097
rect -1461 -1101 -1457 -1097
rect -1454 -1101 -1450 -1097
rect -1447 -1101 -1443 -1097
rect -1440 -1101 -1436 -1097
rect -1433 -1101 -1429 -1097
rect -1496 -1225 -1492 -1221
rect -1475 -1225 -1471 -1221
rect -1468 -1225 -1464 -1221
rect -1461 -1225 -1457 -1221
rect -1454 -1225 -1450 -1221
rect -1447 -1225 -1443 -1221
rect -1440 -1225 -1436 -1221
rect -1433 -1225 -1429 -1221
rect -2408 -1460 -2313 -1331
rect -1817 -1401 -1679 -1388
rect -1683 -1403 -1679 -1401
rect -427 -1453 -419 -1451
rect -427 -1454 -425 -1453
rect -527 -1475 -524 -1460
rect -458 -1464 -454 -1461
rect -414 -1475 -411 -1445
rect -527 -1478 -411 -1475
rect -397 -1496 -392 -145
rect -1393 -1501 -392 -1496
rect -1393 -1817 -1380 -1501
rect -384 -1504 -379 -137
rect -1084 -1509 -379 -1504
rect -1393 -1819 -1381 -1817
rect -1084 -1820 -1071 -1509
rect -371 -1512 -366 -129
rect -775 -1517 -366 -1512
rect -775 -1819 -762 -1517
rect -358 -1520 -353 -121
rect -345 -1496 -340 -113
rect -332 -1365 -327 -100
rect -332 -1374 -327 -1369
rect -319 -148 -314 -87
rect 58 -95 63 1248
rect 80 1245 83 1304
rect 98 1252 102 1294
rect 176 1255 179 1262
rect 183 1253 186 1304
rect 203 1292 233 1296
rect 229 1167 233 1292
rect 262 1256 266 1296
rect 280 1245 283 1304
rect 376 1255 379 1262
rect 345 1251 349 1254
rect 352 1251 356 1254
rect 359 1251 363 1254
rect 366 1251 370 1254
rect 383 1253 386 1304
rect 492 1261 497 1304
rect 492 1255 496 1261
rect 503 1251 508 1293
rect 535 1293 543 1297
rect 535 1255 539 1293
rect 542 1255 546 1263
rect 758 1229 810 1233
rect 390 1223 394 1226
rect 831 1221 835 1304
rect 382 1195 386 1198
rect 1019 1185 1023 1188
rect 314 1167 318 1178
rect 382 1161 386 1164
rect 758 1105 810 1109
rect 758 981 810 985
rect 758 857 810 861
rect 758 733 810 737
rect 758 609 810 613
rect 758 485 810 489
rect 758 361 810 365
rect 758 237 810 241
rect 1028 229 1029 232
rect 758 113 810 117
rect -319 -1485 -314 -152
rect -306 -100 63 -95
rect 1648 -94 1652 1490
rect 1787 1196 1791 1387
rect 1776 1072 1780 1078
rect -306 -1467 -301 -100
rect 1572 -121 1621 -117
rect 1572 -148 1576 -121
rect 1588 -134 1629 -130
rect 1588 -184 1591 -134
rect 1607 -173 1646 -169
rect 1519 -188 1595 -184
rect 1519 -221 1522 -188
rect 1607 -211 1654 -208
rect -273 -223 -269 -222
rect 1650 -222 1654 -211
rect 1686 -222 1690 -173
rect 1706 -353 1710 200
rect 1706 -1072 1710 -357
rect 1706 -1349 1710 -1085
rect 1716 -477 1720 324
rect 1716 -763 1720 -481
rect 1716 -1349 1720 -776
rect 1726 -454 1730 448
rect 1726 -601 1730 -467
rect 1726 -1349 1730 -605
rect 1736 -145 1740 572
rect 1736 -725 1740 -158
rect 1736 -1349 1740 -729
rect 1746 164 1750 696
rect 1746 -849 1750 151
rect 1746 -1349 1750 -853
rect 1757 473 1761 820
rect 1757 -973 1761 460
rect 1757 -1349 1761 -977
rect 1767 782 1771 944
rect 1767 -1097 1771 769
rect 1767 -1349 1771 -1101
rect 1776 -1221 1780 1068
rect 1776 -1349 1780 -1225
rect 1787 -1345 1791 1192
rect 1796 80 1800 1320
rect 2318 1316 2449 1462
rect 2318 1021 2449 1167
rect 2330 718 2461 864
rect 2351 404 2482 550
rect 2325 90 2456 236
rect 1796 -229 1800 76
rect 2334 -200 2465 -54
rect 1796 -1381 1800 -233
rect 2327 -529 2458 -383
rect 2323 -838 2454 -692
rect 2308 -1138 2439 -992
rect 1796 -1394 1817 -1381
rect 1528 -1454 1532 -1450
rect 1535 -1454 1539 -1450
rect 1542 -1454 1546 -1450
rect 1549 -1454 1553 -1450
rect 1618 -1454 1621 -1450
rect 1519 -1467 1522 -1460
rect 1580 -1485 1584 -1462
rect 1588 -1492 1592 -1462
rect 1643 -1467 1647 -1462
rect 2297 -1464 2428 -1318
rect -345 -1501 -144 -1496
rect -466 -1525 -353 -1520
rect -466 -1817 -453 -1525
rect -157 -1818 -144 -1501
rect 461 -1506 1592 -1492
rect 152 -1820 165 -1546
rect 461 -1817 473 -1506
rect -1467 -2423 -1354 -2322
rect -1135 -2425 -1022 -2324
rect -819 -2404 -706 -2303
rect -524 -2408 -411 -2307
rect -203 -2415 -90 -2314
rect 101 -2409 214 -2308
rect 429 -2409 542 -2308
<< m2contact >>
rect -1395 1446 -1382 1453
rect -473 1386 -460 1393
rect -781 1358 -770 1363
rect -1117 1340 -1059 1355
rect 33 1363 37 1367
rect 199 1350 203 1354
rect 209 1387 213 1391
rect 43 1345 47 1349
rect 207 1328 215 1336
rect 262 1470 266 1474
rect 445 1465 449 1469
rect 454 1440 467 1447
rect 1648 1490 1652 1494
rect 1019 1472 1023 1476
rect 810 1457 817 1461
rect 980 1444 984 1448
rect 763 1426 776 1433
rect 988 1407 992 1411
rect 1071 1407 1075 1411
rect 410 1387 414 1391
rect 1036 1377 1040 1381
rect 1075 1377 1079 1381
rect 1103 1377 1107 1381
rect 425 1350 429 1354
rect 465 1332 469 1336
rect 262 1326 266 1330
rect 543 1344 547 1348
rect 504 1332 508 1336
rect -1638 163 -1634 186
rect -1509 1261 -1504 1266
rect -1564 -84 -1560 -80
rect -1281 1262 -1277 1266
rect -1266 1253 -1262 1257
rect -1144 1262 -1139 1266
rect -984 1262 -979 1266
rect -928 1262 -923 1266
rect -768 1262 -763 1266
rect -517 1294 -513 1298
rect -440 1262 -435 1266
rect 58 1248 63 1252
rect -1496 1139 -1492 1143
rect -1489 1015 -1485 1019
rect -1482 891 -1478 895
rect -1475 767 -1471 771
rect -1468 643 -1464 647
rect -1461 519 -1457 523
rect -1454 395 -1450 399
rect -1447 271 -1443 275
rect -1440 147 -1436 151
rect -1433 23 -1429 27
rect -1533 -111 -1529 -107
rect -484 1171 -478 1175
rect -497 1163 -491 1167
rect -1637 -170 -1633 -166
rect -527 -222 -523 -218
rect -1516 -226 -1512 -222
rect -1424 -226 -1420 -222
rect -1433 -233 -1429 -229
rect -1761 -291 -1757 -287
rect -1566 -343 -1562 -339
rect -1440 -357 -1436 -353
rect -1768 -415 -1764 -411
rect -1447 -481 -1443 -477
rect -1775 -539 -1771 -535
rect -1454 -605 -1450 -601
rect -1782 -663 -1778 -659
rect -1461 -729 -1457 -725
rect -1789 -787 -1785 -783
rect -1468 -853 -1464 -849
rect -1796 -911 -1792 -907
rect -1475 -977 -1471 -973
rect -1803 -1035 -1799 -1031
rect -1482 -1101 -1478 -1097
rect -1810 -1159 -1806 -1155
rect -1489 -1225 -1485 -1221
rect -1817 -1283 -1813 -1279
rect -1496 -1349 -1492 -1345
rect -1683 -1407 -1679 -1403
rect -416 -1445 -411 -1440
rect -1626 -1463 -1622 -1457
rect -466 -1466 -462 -1462
rect -425 -1459 -419 -1453
rect -458 -1468 -454 -1464
rect -332 -1369 -327 -1365
rect 98 1294 102 1298
rect 175 1262 180 1266
rect 106 1256 110 1260
rect 262 1296 266 1300
rect 199 1292 203 1296
rect 262 1252 266 1256
rect 375 1262 380 1266
rect 306 1256 310 1260
rect 504 1293 508 1297
rect 543 1293 547 1297
rect 542 1263 546 1267
rect 806 1238 810 1242
rect 754 1229 758 1233
rect 229 1163 233 1167
rect 314 1163 318 1167
rect 806 1114 810 1118
rect 754 1105 758 1109
rect 806 990 810 994
rect 754 981 758 985
rect 806 866 810 870
rect 754 857 758 861
rect 806 742 810 746
rect 754 733 758 737
rect 806 618 810 622
rect 754 609 758 613
rect 806 494 810 498
rect 754 485 758 489
rect 806 370 810 374
rect 754 361 758 365
rect 806 246 810 250
rect 754 237 758 241
rect 806 122 810 126
rect 754 113 758 117
rect -319 -152 -314 -148
rect 1787 1387 1791 1400
rect 1813 1387 1818 1400
rect 1787 1192 1791 1196
rect 1776 1078 1780 1091
rect 1776 1068 1780 1072
rect 1767 944 1771 948
rect 1757 820 1761 824
rect 1746 696 1750 700
rect 1736 572 1740 576
rect 1726 448 1730 452
rect 1716 324 1720 328
rect 1706 200 1710 204
rect 1572 -152 1576 -148
rect 1694 -159 1698 -155
rect -273 -222 -269 -218
rect 1693 -222 1697 -218
rect 1706 -357 1710 -353
rect 1706 -1085 1710 -1072
rect 1716 -481 1720 -477
rect 1716 -776 1720 -763
rect 1726 -467 1730 -454
rect 1726 -605 1730 -601
rect 1736 -158 1740 -145
rect 1736 -729 1740 -725
rect 1746 151 1750 164
rect 1746 -853 1750 -849
rect 1757 460 1761 473
rect 1757 -977 1761 -973
rect 1767 769 1771 782
rect 1767 -1101 1771 -1097
rect 1776 -1225 1780 -1221
rect 1787 -1349 1791 -1345
rect 1813 1078 1817 1091
rect 1813 769 1817 782
rect 1813 460 1817 473
rect 1813 151 1817 164
rect 1796 76 1800 80
rect 1813 -158 1817 -145
rect 1796 -233 1800 -229
rect 1813 -467 1817 -454
rect 1813 -776 1817 -763
rect 1813 -1085 1817 -1072
rect 1643 -1444 1647 -1440
rect 1693 -1444 1697 -1440
rect 1572 -1455 1576 -1451
rect 1621 -1454 1625 -1450
rect -306 -1472 -301 -1467
rect 1519 -1472 1524 -1467
rect -319 -1489 -314 -1485
rect 1580 -1489 1584 -1485
rect 1643 -1472 1647 -1467
rect 152 -1546 165 -1538
<< metal2 >>
rect -1509 1275 -1484 1909
rect -50 1453 -47 1504
rect -1382 1446 -47 1453
rect -34 1433 -31 1504
rect -18 1447 -15 1504
rect -2 1486 1 1496
rect 14 1493 17 1496
rect 239 1493 242 1499
rect 14 1490 242 1493
rect 247 1486 250 1499
rect -2 1483 250 1486
rect 255 1460 258 1499
rect 263 1474 266 1499
rect 271 1468 274 1499
rect 279 1476 282 1499
rect 287 1494 290 1499
rect 295 1494 298 1499
rect 295 1490 1648 1494
rect 279 1473 1019 1476
rect 271 1465 445 1468
rect 255 1457 810 1460
rect -18 1440 454 1447
rect -34 1426 763 1433
rect 59 1387 209 1391
rect 37 1363 183 1367
rect -1116 1275 -1059 1340
rect -513 1294 98 1298
rect 199 1296 203 1350
rect 207 1275 215 1328
rect 262 1300 266 1326
rect 425 1275 429 1350
rect 469 1332 504 1336
rect 504 1297 508 1332
rect 535 1275 539 1332
rect 543 1297 547 1344
rect 988 1275 992 1407
rect 1075 1407 1087 1411
rect 1071 1389 1075 1407
rect 1061 1385 1075 1389
rect 1791 1387 1813 1400
rect 1061 1381 1065 1385
rect 1040 1377 1065 1381
rect 1079 1377 1103 1381
rect -1509 1267 992 1275
rect -1509 1266 542 1267
rect -1504 1262 -1281 1266
rect -1277 1262 -1144 1266
rect -1139 1262 -984 1266
rect -979 1262 -928 1266
rect -923 1262 -768 1266
rect -763 1262 -440 1266
rect -435 1262 175 1266
rect 180 1262 375 1266
rect 380 1263 542 1266
rect 546 1263 992 1267
rect 380 1262 992 1263
rect -1504 1261 992 1262
rect 1004 1312 1036 1316
rect -1386 1238 -1382 1261
rect -1386 1234 -1378 1238
rect -1244 1234 -1240 1261
rect -1085 1234 -1081 1261
rect -868 1234 -864 1261
rect -541 1234 -537 1261
rect 74 1234 78 1261
rect 106 1260 110 1261
rect 274 1234 278 1261
rect 306 1260 310 1261
rect 430 1188 491 1192
rect 226 1163 229 1167
rect 233 1163 314 1167
rect -1492 1139 -1378 1143
rect -1234 1139 -1230 1143
rect -1214 1139 -1208 1143
rect -1069 1138 -1062 1143
rect -1054 1139 -1048 1143
rect -859 1139 -852 1144
rect 23 1143 30 1144
rect -534 1138 -527 1143
rect 14 1139 82 1143
rect 214 1140 252 1143
rect 430 1143 435 1188
rect 754 1143 758 1229
rect 258 1140 282 1143
rect 214 1139 282 1140
rect 414 1139 758 1143
rect 770 1142 773 1261
rect 1004 1252 1008 1312
rect 805 1238 806 1242
rect 1151 1192 1787 1196
rect 770 1139 823 1142
rect 805 1114 806 1118
rect 430 1064 490 1068
rect -1485 1015 -1378 1019
rect -1214 1015 -1208 1019
rect -1054 1015 -1048 1019
rect 14 1015 82 1019
rect 214 1016 252 1019
rect 430 1019 435 1064
rect 754 1019 758 1105
rect 1780 1078 1813 1091
rect 1151 1068 1776 1072
rect 258 1016 282 1019
rect 214 1015 282 1016
rect 412 1015 758 1019
rect 805 990 806 994
rect 430 940 490 944
rect -1478 891 -1371 895
rect -1214 891 -1208 895
rect -1054 891 -1048 895
rect 14 891 82 895
rect 214 892 252 895
rect 430 895 435 940
rect 754 895 758 981
rect 1151 944 1767 948
rect 258 892 282 895
rect 214 891 282 892
rect 412 891 758 895
rect 805 866 806 870
rect 430 816 490 820
rect -1471 767 -1364 771
rect -1214 767 -1208 771
rect -1054 767 -1048 771
rect 14 767 82 771
rect 214 768 252 771
rect 430 771 435 816
rect 754 771 758 857
rect 1151 820 1757 824
rect 258 768 282 771
rect 214 767 282 768
rect 412 767 758 771
rect 1771 769 1813 782
rect 805 742 806 746
rect 430 692 490 696
rect -1464 643 -1357 647
rect -1214 643 -1208 647
rect -1054 643 -1048 647
rect 14 643 82 647
rect 214 644 252 647
rect 430 647 435 692
rect 754 647 758 733
rect 1151 696 1746 700
rect 258 644 282 647
rect 214 643 282 644
rect 412 643 758 647
rect 805 618 806 622
rect 430 568 490 572
rect -1457 519 -1350 523
rect -1214 519 -1208 523
rect -1054 519 -1048 523
rect 14 519 82 523
rect 214 520 252 523
rect 430 523 435 568
rect 754 523 758 609
rect 1151 572 1736 576
rect 258 520 282 523
rect 214 519 282 520
rect 412 519 758 523
rect 805 494 806 498
rect 430 444 490 448
rect -1450 395 -1343 399
rect -1214 395 -1208 399
rect -1054 395 -1048 399
rect 14 395 82 399
rect 214 396 252 399
rect 430 399 435 444
rect 754 399 758 485
rect 1761 460 1813 473
rect 1151 448 1726 452
rect 258 396 282 399
rect 214 395 282 396
rect 412 395 758 399
rect 805 370 806 374
rect 430 320 490 324
rect -1443 271 -1336 275
rect -1214 271 -1208 275
rect -1054 271 -1048 275
rect 14 271 82 275
rect 214 272 252 275
rect 430 275 435 320
rect 754 275 758 361
rect 1151 324 1716 328
rect 258 272 282 275
rect 214 271 282 272
rect 412 271 758 275
rect 805 246 806 250
rect 430 196 490 200
rect -1942 163 -1638 186
rect -1436 147 -1329 151
rect -1214 147 -1208 151
rect -1054 147 -1048 151
rect 14 147 82 151
rect 214 148 252 151
rect 430 151 435 196
rect 754 151 758 237
rect 1151 200 1706 204
rect 1750 151 1813 164
rect 258 148 282 151
rect 214 147 282 148
rect 412 147 758 151
rect 805 122 806 126
rect 430 72 490 76
rect -1429 23 -1322 27
rect -1214 23 -1208 27
rect -1054 23 -1048 27
rect 14 23 82 27
rect 214 24 252 27
rect 430 27 435 72
rect 754 27 758 113
rect 1151 76 1796 80
rect 1800 76 1805 80
rect 258 24 282 27
rect 214 23 282 24
rect 412 23 758 27
rect 1007 13 1010 23
rect -1533 -152 -1529 -111
rect 1615 -151 1653 -147
rect -1633 -170 -1544 -166
rect 1615 -176 1619 -151
rect 1740 -158 1813 -145
rect -523 -222 -273 -218
rect 1505 -221 1508 -203
rect 1694 -218 1697 -159
rect -1512 -226 -1424 -222
rect -1496 -233 -1433 -229
rect -1429 -233 -1425 -229
rect -426 -233 -275 -229
rect 1556 -283 1560 -229
rect 1653 -233 1796 -229
rect 1699 -283 1703 -233
rect -1757 -291 -1568 -287
rect -1562 -343 -1415 -340
rect -523 -343 -214 -340
rect -1496 -357 -1440 -353
rect -1436 -357 -1425 -353
rect -426 -357 -275 -353
rect 1554 -357 1565 -353
rect 1654 -357 1706 -353
rect 1710 -357 1716 -353
rect 1556 -407 1560 -357
rect 1699 -407 1703 -357
rect -1764 -415 -1568 -411
rect -530 -467 -197 -464
rect 1730 -467 1813 -454
rect -1496 -481 -1447 -477
rect -1443 -481 -1425 -477
rect -426 -481 -275 -477
rect 1554 -481 1565 -477
rect 1638 -481 1716 -477
rect 1720 -481 1726 -477
rect 1556 -531 1560 -481
rect 1699 -531 1703 -481
rect -1771 -539 -1568 -535
rect -530 -591 -197 -588
rect -1496 -605 -1454 -601
rect -1450 -605 -1425 -601
rect -426 -605 -275 -601
rect 1554 -605 1565 -601
rect 1638 -605 1726 -601
rect 1730 -605 1736 -601
rect 1556 -655 1560 -605
rect 1699 -655 1703 -605
rect -1778 -663 -1568 -659
rect -530 -715 -197 -712
rect -1496 -729 -1461 -725
rect -1457 -729 -1425 -725
rect -426 -729 -275 -725
rect 1554 -729 1565 -725
rect 1629 -729 1736 -725
rect 1740 -729 1746 -725
rect 1556 -779 1560 -729
rect 1699 -779 1703 -729
rect 1720 -776 1813 -763
rect -1785 -787 -1568 -783
rect -530 -839 -197 -836
rect -1496 -853 -1468 -849
rect -1464 -853 -1425 -849
rect -426 -853 -275 -849
rect 1554 -853 1565 -849
rect 1634 -853 1746 -849
rect 1750 -853 1757 -849
rect 1556 -903 1560 -853
rect 1699 -903 1703 -853
rect -1792 -911 -1568 -907
rect -530 -963 -197 -960
rect -1496 -977 -1475 -973
rect -1471 -977 -1425 -973
rect -426 -977 -275 -973
rect 1554 -977 1565 -973
rect 1631 -977 1757 -973
rect 1761 -977 1767 -973
rect 1556 -1027 1560 -977
rect 1699 -1027 1703 -977
rect -1799 -1035 -1568 -1031
rect -530 -1087 -197 -1084
rect 1710 -1085 1813 -1072
rect -1496 -1101 -1482 -1097
rect -1478 -1101 -1425 -1097
rect -426 -1101 -275 -1097
rect 1554 -1101 1565 -1097
rect 1624 -1101 1767 -1097
rect 1771 -1101 1776 -1097
rect 1556 -1151 1560 -1101
rect 1699 -1151 1703 -1101
rect -1806 -1159 -1568 -1155
rect -530 -1211 -197 -1208
rect -1496 -1225 -1489 -1221
rect -1485 -1225 -1425 -1221
rect -426 -1225 -275 -1221
rect 1554 -1225 1565 -1221
rect 1628 -1225 1776 -1221
rect 1780 -1225 1787 -1221
rect 1556 -1275 1560 -1225
rect 1699 -1275 1703 -1225
rect -1813 -1283 -1568 -1279
rect -530 -1335 -197 -1332
rect -1492 -1349 -1425 -1345
rect -426 -1349 -275 -1345
rect 1625 -1349 1787 -1345
rect 1791 -1349 1796 -1345
rect 1556 -1381 1560 -1349
rect 1699 -1399 1703 -1349
rect -1679 -1407 -1568 -1403
rect -426 -1444 -416 -1440
rect 1620 -1444 1643 -1440
rect 1668 -1444 1693 -1440
rect 1668 -1450 1671 -1444
rect 1618 -1454 1621 -1450
rect 1625 -1454 1671 -1450
rect 1572 -1456 1576 -1455
rect -419 -1459 -197 -1456
rect 1522 -1460 1576 -1456
rect -466 -1489 -462 -1466
rect -458 -1472 -418 -1468
rect 1524 -1472 1643 -1467
rect -423 -1538 -418 -1472
rect -423 -1545 152 -1538
rect -117 -1546 152 -1545
<< m3contact >>
rect 286 1490 290 1494
rect 976 1444 980 1448
rect 406 1387 410 1391
rect -473 1382 -460 1386
rect -781 1353 -770 1358
rect 43 1341 47 1345
rect 58 1252 63 1256
rect 258 1252 262 1256
rect -484 1175 -478 1179
rect 222 1163 226 1167
rect 252 1140 258 1146
rect 801 1238 805 1242
rect 801 1114 805 1118
rect 252 1016 258 1022
rect 801 990 805 994
rect 252 892 258 898
rect 801 866 805 870
rect 252 768 258 774
rect 801 742 805 746
rect 252 644 258 650
rect 801 618 805 622
rect 252 520 258 526
rect 801 494 805 498
rect 252 396 258 402
rect 801 370 805 374
rect 252 272 258 278
rect 801 246 805 250
rect -1956 163 -1942 186
rect 252 148 258 154
rect 801 122 805 126
rect 252 24 258 30
rect -1564 -80 -1560 -76
rect -1533 -156 -1529 -152
rect -819 -156 -814 -152
rect -319 -156 -314 -152
rect 1572 -156 1576 -152
rect 1556 -287 1560 -283
rect 1556 -411 1560 -407
rect 1556 -535 1560 -531
rect 1556 -659 1560 -655
rect 1556 -783 1560 -779
rect 1556 -907 1560 -903
rect 1556 -1031 1560 -1027
rect 1556 -1155 1560 -1151
rect 1556 -1279 1560 -1275
rect -332 -1373 -327 -1369
rect 1556 -1385 1560 -1381
rect -1622 -1462 -1618 -1458
rect -306 -1467 -301 -1463
rect -466 -1493 -462 -1489
rect -319 -1493 -314 -1489
rect 1580 -1493 1584 -1489
<< metal3 >>
rect -1565 1494 291 1495
rect -1565 1490 286 1494
rect 290 1490 291 1494
rect -1565 1489 291 1490
rect -1957 186 -1941 187
rect -1957 163 -1956 186
rect -1942 163 -1941 186
rect -1957 162 -1941 163
rect -1565 -76 -1559 1489
rect 975 1448 981 1449
rect 975 1444 976 1448
rect 980 1444 981 1448
rect 975 1392 981 1444
rect 313 1391 981 1392
rect 313 1387 406 1391
rect 410 1387 981 1391
rect -1401 1386 -459 1387
rect -1401 1382 -473 1386
rect -460 1382 -459 1386
rect -1401 1381 -459 1382
rect 313 1386 981 1387
rect -1401 1168 -1395 1381
rect -782 1358 -769 1359
rect -782 1353 -781 1358
rect -770 1353 -769 1358
rect -782 1288 -769 1353
rect 42 1345 48 1346
rect 42 1341 43 1345
rect 47 1341 48 1345
rect 42 1288 48 1341
rect 313 1288 319 1386
rect -1343 1282 319 1288
rect -1367 1251 -520 1257
rect -485 1179 -477 1282
rect 57 1256 294 1257
rect 57 1252 58 1256
rect 63 1252 258 1256
rect 262 1252 294 1256
rect 57 1251 294 1252
rect -485 1175 -484 1179
rect -478 1175 -477 1179
rect -485 1174 -477 1175
rect 251 1242 806 1243
rect 251 1238 801 1242
rect 805 1238 806 1242
rect 251 1237 806 1238
rect -1401 1167 227 1168
rect -1401 1163 222 1167
rect 226 1163 227 1167
rect -1401 1162 227 1163
rect 251 1146 259 1237
rect 251 1140 252 1146
rect 258 1140 259 1146
rect 251 1139 259 1140
rect 251 1118 806 1119
rect 251 1114 801 1118
rect 805 1114 806 1118
rect 251 1113 806 1114
rect 251 1022 259 1113
rect 251 1016 252 1022
rect 258 1016 259 1022
rect 251 1015 259 1016
rect 251 994 806 995
rect 251 990 801 994
rect 805 990 806 994
rect 251 989 806 990
rect 251 898 259 989
rect 251 892 252 898
rect 258 892 259 898
rect 251 891 259 892
rect 251 870 806 871
rect 251 866 801 870
rect 805 866 806 870
rect 251 865 806 866
rect 251 774 259 865
rect 251 768 252 774
rect 258 768 259 774
rect 251 767 259 768
rect 251 746 806 747
rect 251 742 801 746
rect 805 742 806 746
rect 251 741 806 742
rect 251 650 259 741
rect 251 644 252 650
rect 258 644 259 650
rect 251 643 259 644
rect 251 622 806 623
rect 251 618 801 622
rect 805 618 806 622
rect 251 617 806 618
rect 251 526 259 617
rect 251 520 252 526
rect 258 520 259 526
rect 251 519 259 520
rect 251 498 806 499
rect 251 494 801 498
rect 805 494 806 498
rect 251 493 806 494
rect 251 402 259 493
rect 251 396 252 402
rect 258 396 259 402
rect 251 395 259 396
rect 251 374 806 375
rect 251 370 801 374
rect 805 370 806 374
rect 251 369 806 370
rect 251 278 259 369
rect 251 272 252 278
rect 258 272 259 278
rect 251 271 259 272
rect 251 250 806 251
rect 251 246 801 250
rect 805 246 806 250
rect 251 245 806 246
rect 251 154 259 245
rect 251 148 252 154
rect 258 148 259 154
rect 251 147 259 148
rect 251 126 806 127
rect 251 122 801 126
rect 805 122 806 126
rect 251 121 806 122
rect 251 30 259 121
rect 595 75 602 81
rect 251 24 252 30
rect 258 24 259 30
rect 251 23 259 24
rect -1565 -80 -1564 -76
rect -1560 -80 -1559 -76
rect -1565 -81 -1559 -80
rect -1534 -152 1577 -151
rect -1534 -156 -1533 -152
rect -1529 -156 -819 -152
rect -814 -156 -319 -152
rect -314 -156 1572 -152
rect 1576 -156 1577 -152
rect -1534 -157 1577 -156
rect 1555 -283 1561 -282
rect -1505 -287 1556 -283
rect 1560 -287 1640 -283
rect -1505 -288 1640 -287
rect 1555 -407 1561 -406
rect -1505 -411 1556 -407
rect 1560 -411 1640 -407
rect -1505 -412 1640 -411
rect 1555 -531 1561 -530
rect 1638 -531 1640 -530
rect -1505 -535 1556 -531
rect 1560 -535 1640 -531
rect -1505 -536 1640 -535
rect 1555 -655 1561 -654
rect 1615 -655 1640 -654
rect -1505 -659 1556 -655
rect 1560 -659 1640 -655
rect -1505 -660 1640 -659
rect 1555 -779 1561 -778
rect 1629 -779 1640 -778
rect -1505 -783 1556 -779
rect 1560 -783 1640 -779
rect -1505 -784 1640 -783
rect 1555 -903 1561 -902
rect 1634 -903 1640 -902
rect -1505 -907 1556 -903
rect 1560 -907 1640 -903
rect -1505 -908 1640 -907
rect 1555 -1027 1561 -1026
rect 1615 -1027 1640 -1026
rect -1505 -1031 1556 -1027
rect 1560 -1031 1640 -1027
rect -1505 -1032 1640 -1031
rect 1555 -1151 1561 -1150
rect 1624 -1151 1640 -1150
rect -1505 -1155 1556 -1151
rect 1560 -1155 1640 -1151
rect -1505 -1156 1640 -1155
rect 1555 -1275 1561 -1274
rect 1628 -1275 1640 -1274
rect -1505 -1279 1556 -1275
rect 1560 -1279 1640 -1275
rect -1505 -1280 1640 -1279
rect -467 -1369 1585 -1368
rect -467 -1373 -332 -1369
rect -327 -1373 1585 -1369
rect -467 -1374 1585 -1373
rect 1555 -1381 1561 -1379
rect 1555 -1385 1556 -1381
rect 1560 -1385 1561 -1381
rect 1555 -1386 1561 -1385
rect 1555 -1399 1560 -1386
rect 1615 -1399 1640 -1398
rect -1505 -1404 1640 -1399
rect -1626 -1458 1609 -1457
rect -1626 -1462 -1622 -1458
rect -1618 -1462 1609 -1458
rect -1626 -1463 1609 -1462
rect -307 -1467 -306 -1463
rect -301 -1467 -300 -1463
rect -307 -1468 -300 -1467
rect -467 -1489 1585 -1488
rect -467 -1493 -466 -1489
rect -462 -1493 -319 -1489
rect -314 -1493 1580 -1489
rect 1584 -1493 1585 -1489
rect -467 -1494 1585 -1493
use inpad  inpad_0
timestamp 1509371954
transform 1 0 -1519 0 1 2183
box -32 -366 277 317
use GNDPad  t1
timestamp 1509371954
transform 1 0 -1242 0 1 1852
box 0 -35 309 648
use InPad  t2
timestamp 1509371954
transform 1 0 -901 0 1 2183
box -32 -366 277 317
use InPad  t3
timestamp 1509371954
transform 1 0 -592 0 1 2183
box -32 -366 277 317
use VddPad  t4
timestamp 1509371954
transform 1 0 -315 0 1 1852
box 0 -35 309 648
use BlankPad  t5
timestamp 1006127261
transform 1 0 5 0 1 1868
box -11 -51 298 632
use inpad  inpad_1
timestamp 1509371954
transform 1 0 335 0 1 2183
box -32 -366 277 317
use inpad  inpad_2
timestamp 1509371954
transform 1 0 644 0 1 2183
box -32 -366 277 317
use outpad  outpad_1
timestamp 1012172318
transform 1 0 904 0 1 1843
box 17 -26 326 657
use outpad  outpad_0
timestamp 1012172318
transform 1 0 1213 0 1 1843
box 17 -26 326 657
use Corner  clt
timestamp 1012241868
transform 1 0 -2325 0 1 1869
box -143 -333 774 618
use fsm  fsm_0
timestamp 1512683710
transform 1 0 -92 0 1 1780
box 0 -285 412 33
use Corner  crt
timestamp 1012241868
transform 0 1 1869 -1 0 2325
box -143 -333 774 618
use inv  inv_0
timestamp 1512712928
transform 0 -1 60 1 0 1392
box -32 -27 3 9
use inv  inv_1
timestamp 1512712928
transform 0 -1 168 1 0 1392
box -32 -27 3 9
use andstat  andstat_0
timestamp 1512636464
transform 1 0 434 0 1 1344
box -12 -14 63 66
use andstat  andstat_1
timestamp 1512636464
transform 1 0 1008 0 1 1401
box -12 -14 63 66
use inv  inv_3
timestamp 1512712928
transform 1 0 1116 0 1 1413
box -32 -27 3 9
use inv  inv_2
timestamp 1512712928
transform 1 0 540 0 1 1355
box -32 -27 3 9
use andstat  andstat_3
timestamp 1512636464
transform -1 0 -1549 0 1 -155
box -12 -14 63 66
use inv  inv_5
timestamp 1512712928
transform 0 1 -1525 -1 0 -195
box -32 -27 3 9
use new_latch  new_latch_3
array 0 0 66 0 9 124
timestamp 1512685536
transform 1 0 -1600 0 1 -1436
box 31 -28 97 96
use bus_10  bus_10_1
timestamp 1512385298
transform 1 0 -1487 0 1 -3407
box -9 1974 58 4676
use phi0_connection  phi0_connection_0
timestamp 1512513482
transform 1 0 -1342 0 1 1265
box -1 -13 5 23
use phi0_connection  phi0_connection_1
timestamp 1512513482
transform 1 0 -1205 0 1 1265
box -1 -13 5 23
use phi0_connection  phi0_connection_2
timestamp 1512513482
transform 1 0 -1045 0 1 1265
box -1 -13 5 23
use phi0_connection  phi0_connection_3
timestamp 1512513482
transform 1 0 -829 0 1 1265
box -1 -13 5 23
use phi0_connection  phi0_connection_4
timestamp 1512513482
transform 1 0 -501 0 1 1265
box -1 -13 5 23
use phi1_connection  phi1_connection_4
timestamp 1512512927
transform 1 0 -1346 0 1 1169
box 3 -7 9 13
use phi1_connection  phi1_connection_5
timestamp 1512512927
transform 1 0 -1209 0 1 1169
box 3 -7 9 13
use phi1_connection  phi1_connection_3
timestamp 1512512927
transform 1 0 -1049 0 1 1169
box 3 -7 9 13
use phi1_connection  phi1_connection_2
timestamp 1512512927
transform 1 0 -833 0 1 1169
box 3 -7 9 13
use phi1_connection  phi1_connection_1
timestamp 1512512927
transform 1 0 -505 0 1 1169
box 3 -7 9 13
use sreg_01  sreg_01_0
timestamp 1512534937
transform 1 0 -1283 0 1 12
box -95 3 42 1247
use sreg_02  sreg_02_0
timestamp 1512534937
transform 1 0 -1146 0 1 12
box -95 0 65 1248
use sreg_04  sreg_04_0
timestamp 1512539734
transform 1 0 -986 0 1 12
box -95 0 121 1248
use sreg_08  sreg_08_0
timestamp 1512534937
transform 1 0 -770 0 1 12
box -95 0 233 1248
use sreg_16  sreg_16_0
timestamp 1512534937
transform 1 0 -442 0 1 12
box -95 0 457 1248
use phi0_connection  phi0_connection_5
timestamp 1512513482
transform 1 0 114 0 1 1265
box -1 -13 5 23
use phi1_connection  phi1_connection_0
timestamp 1512512927
transform 1 0 110 0 1 1169
box 3 -7 9 13
use sreg_01  sreg_01_1
timestamp 1512534937
transform 1 0 173 0 1 12
box -95 3 42 1247
use phi0_connection  phi0_connection_6
timestamp 1512513482
transform 1 0 314 0 1 1265
box -1 -13 5 23
use sreg_01  sreg_01_2
timestamp 1512534937
transform 1 0 373 0 1 12
box -95 3 42 1247
use sreg_out_connection  sreg_out_connection_9
timestamp 1512685257
transform 1 0 587 0 1 1175
box -38 16 565 22
use add_latch_connections  add_latch_connections_9
timestamp 1512633651
transform 1 0 1009 0 1 1222
box -1 -83 81 2
use sreg_out_connection  sreg_out_connection_0
timestamp 1512685257
transform 1 0 587 0 1 1051
box -38 16 565 22
use add_latch_connections  add_latch_connections_8
timestamp 1512633651
transform 1 0 1009 0 1 1098
box -1 -83 81 2
use sreg_out_connection  sreg_out_connection_1
timestamp 1512685257
transform 1 0 587 0 1 927
box -38 16 565 22
use add_latch_connections  add_latch_connections_7
timestamp 1512633651
transform 1 0 1009 0 1 974
box -1 -83 81 2
use sreg_out_connection  sreg_out_connection_2
timestamp 1512685257
transform 1 0 587 0 1 803
box -38 16 565 22
use add_latch_connections  add_latch_connections_6
timestamp 1512633651
transform 1 0 1009 0 1 850
box -1 -83 81 2
use sreg_out_connection  sreg_out_connection_3
timestamp 1512685257
transform 1 0 587 0 1 679
box -38 16 565 22
use add_latch_connections  add_latch_connections_5
timestamp 1512633651
transform 1 0 1009 0 1 726
box -1 -83 81 2
use sreg_out_connection  sreg_out_connection_4
timestamp 1512685257
transform 1 0 587 0 1 555
box -38 16 565 22
use add_latch_connections  add_latch_connections_4
timestamp 1512633651
transform 1 0 1009 0 1 602
box -1 -83 81 2
use sreg_out_connection  sreg_out_connection_5
timestamp 1512685257
transform 1 0 587 0 1 431
box -38 16 565 22
use add_latch_connections  add_latch_connections_3
timestamp 1512633651
transform 1 0 1009 0 1 478
box -1 -83 81 2
use sreg_out_connection  sreg_out_connection_6
timestamp 1512685257
transform 1 0 587 0 1 307
box -38 16 565 22
use add_latch_connections  add_latch_connections_2
timestamp 1512633651
transform 1 0 1009 0 1 354
box -1 -83 81 2
use sreg_out_connection  sreg_out_connection_7
timestamp 1512685257
transform 1 0 587 0 1 183
box -38 16 565 22
use add_latch_connections  add_latch_connections_1
timestamp 1512633651
transform 1 0 1009 0 1 230
box -1 -83 81 2
use sreg_out_connection  sreg_out_connection_8
timestamp 1512685257
transform 1 0 587 0 1 59
box -38 16 565 22
use new_latch  new_latch_0
array 0 0 102 0 9 124
timestamp 1512685536
transform 1 0 458 0 1 43
box 31 -28 97 96
use add_latch_connections  add_latch_connections_0
timestamp 1512633651
transform 1 0 1009 0 1 106
box -1 -83 81 2
use addsub_eight  addsub_eight_0
timestamp 1512379736
transform 1 0 810 0 1 14
box 4 -1 200 1239
use latch_shift  latch_shift_0
array 0 0 66 0 10 124
timestamp 1512686560
transform 1 0 1002 0 -1 1359
box 31 -28 97 163
use andstat  andstat_2
timestamp 1512636464
transform 1 0 1637 0 1 -165
box -12 -14 63 66
use inv  inv_4
timestamp 1512712928
transform 0 1 1618 -1 0 -205
box -32 -27 3 9
use phi1_connection  phi1_connection_6
timestamp 1512512927
transform -1 0 -458 0 -1 -1375
box 3 -7 9 13
use sreg_32  sreg_32_0
timestamp 1512534937
transform -1 0 -521 0 -1 -218
box -95 0 905 1248
use phi1_connection  phi1_connection_7
timestamp 1512512927
transform -1 0 1588 0 -1 -1375
box 3 -7 9 13
use sreg_64  sreg_64_0
timestamp 1512538665
transform -1 0 1525 0 -1 -218
box -95 0 1801 1248
use new_latch  new_latch_2
array 0 0 -66 0 9 -124
timestamp 1512685536
transform -1 0 1731 0 -1 -1366
box 31 -28 97 96
use outPad  outPad_1
array 0 9 -309 0 0 683
timestamp 1012172318
transform 0 1 1843 -1 0 -1213
box 17 -26 326 657
use InPad  InPad_1
array 0 9 309 0 0 -683
timestamp 1509371954
transform 0 -1 -2183 1 0 -1520
box -32 -366 277 317
use Corner  clb
timestamp 1012241868
transform 0 -1 -1869 1 0 -2325
box -143 -333 774 618
use Corner  crb
timestamp 1012241868
transform -1 0 2325 0 -1 -1869
box -143 -333 774 618
use InPad  InPad_2
array 0 9 -309 0 0 -683
timestamp 1509371954
transform -1 0 -1261 0 -1 -2183
box -32 -366 277 317
<< labels >>
rlabel metal1 -460 2372 -460 2372 1 phi1
rlabel metal1 -1428 2373 -1427 2373 1 RESET
rlabel metal1 462 2377 462 2377 1 iter
rlabel metal1 755 2377 755 2377 1 load
rlabel metal1 1066 2371 1066 2372 1 ready
rlabel metal1 -1423 -2394 -1423 -2394 1 bp0
rlabel metal1 -1097 -2388 -1097 -2388 1 bp1
rlabel metal1 -782 -2379 -782 -2379 1 bp2
rlabel metal1 -487 -2360 -487 -2360 1 bp3
rlabel metal1 -156 -2373 -156 -2373 1 bp4
rlabel metal1 146 -2370 146 -2370 1 bp5
rlabel metal1 481 -2368 481 -2368 1 bp6
rlabel metal1 -2372 1385 -2372 1385 1 in0
rlabel metal1 -2374 1079 -2374 1079 1 in1
rlabel metal1 -2365 737 -2365 737 1 in2
rlabel metal1 -2341 435 -2341 435 1 in3
rlabel metal1 -2351 123 -2351 123 1 in4
rlabel metal1 -2362 -205 -2362 -205 1 in5
rlabel metal1 -2379 -493 -2379 -493 1 in6
rlabel metal1 -2386 -819 -2386 -819 1 in7
rlabel metal1 -2367 -1107 -2367 -1107 1 in8
rlabel metal1 -2377 -1405 -2377 -1405 1 in9
rlabel metal1 2367 -1405 2367 -1405 1 out0
rlabel metal1 2365 -1084 2365 -1084 1 out1
rlabel metal1 2388 -784 2388 -784 1 out2
rlabel metal1 2376 -461 2376 -461 1 out3
rlabel metal1 2374 -161 2374 -161 1 out4
rlabel metal1 2381 139 2381 139 1 out5
rlabel metal1 2400 456 2400 456 1 out6
rlabel metal1 2379 765 2379 765 1 out7
rlabel metal1 2369 1070 2369 1070 1 out8
rlabel metal1 2355 1365 2355 1365 1 out9
rlabel metal1 1364 2382 1364 2382 1 out10
rlabel metal1 53 1460 53 1460 1 p2-
rlabel metal1 202 1460 202 1460 1 p1
rlabel metal1 193 1460 193 1460 1 p1-
rlabel metal1 -778 2364 -778 2364 1 phi0
rlabel metal1 265 1467 265 1467 1 sreg_en
rlabel metal2 273 1469 273 1469 1 sreg_latch
rlabel metal2 281 1474 281 1474 1 add_latch
rlabel metal2 -286 -1347 -286 -1347 1 o64_0
rlabel metal3 -1501 -1401 -1501 -1401 1 input_latch_9
rlabel metal1 1551 -1452 1551 -1452 1 64_c0
rlabel metal1 1544 -1452 1544 -1452 1 64_c0-
rlabel metal1 1537 -1452 1537 -1452 1 64_c1
rlabel metal1 1530 -1452 1530 -1452 1 64_c1-
rlabel metal2 -241 -1333 -241 -1333 8 Vdd!_uq0
rlabel metal2 -212 -1333 -212 -1333 8 Vdd!_uq0
rlabel metal2 -522 -1333 -522 -1333 8 Vdd!_uq0
rlabel metal2 -241 -1085 -241 -1085 8 Vdd!_uq1
rlabel metal2 -212 -1085 -212 -1085 8 Vdd!_uq1
rlabel metal2 -522 -1085 -522 -1085 8 Vdd!_uq1
rlabel metal2 -241 -961 -241 -961 8 Vdd!_uq2
rlabel metal2 -212 -961 -212 -961 8 Vdd!_uq2
rlabel metal2 -522 -961 -522 -961 8 Vdd!_uq2
rlabel metal2 -241 -837 -241 -837 8 Vdd!_uq3
rlabel metal2 -212 -837 -212 -837 8 Vdd!_uq3
rlabel metal2 -522 -837 -522 -837 8 Vdd!_uq3
rlabel metal2 -241 -713 -241 -713 8 Vdd!_uq4
rlabel metal2 -212 -713 -212 -713 8 Vdd!_uq4
rlabel metal2 -522 -713 -522 -713 8 Vdd!_uq4
rlabel metal2 -241 -589 -241 -589 8 Vdd!_uq5
rlabel metal2 -212 -589 -212 -589 8 Vdd!_uq5
rlabel metal2 -522 -589 -522 -589 8 Vdd!_uq5
rlabel metal2 -241 -465 -241 -465 8 Vdd!_uq6
rlabel metal2 -212 -465 -212 -465 8 Vdd!_uq6
rlabel metal2 -522 -465 -522 -465 8 Vdd!_uq6
rlabel metal2 -241 -1457 -241 -1457 8 Vdd!_uq8
rlabel metal2 -212 -1457 -212 -1457 8 Vdd!_uq8
rlabel metal1 -1392 1983 -1392 1983 1 in_uq3
rlabel metal1 -779 1983 -779 1983 1 in_uq13
rlabel m2contact -1494 -1347 -1494 -1347 1 32_bit9
rlabel metal2 -1232 1140 -1232 1140 1 1_bit9
rlabel metal2 432 1141 432 1141 1 last_bit9
rlabel metal2 27 1141 27 1141 1 16_bit9
rlabel metal2 -1066 1140 -1065 1140 1 2_bit9
rlabel metal2 -855 1140 -855 1140 1 4_bit9
rlabel metal2 -530 1141 -530 1141 1 8_bit9
rlabel metal1 -1172 1248 -1172 1248 1 2_c0
rlabel metal1 -1165 1248 -1165 1248 1 2_c0-
rlabel metal1 -1158 1248 -1158 1248 1 2_c1
rlabel metal1 -1151 1248 -1151 1248 1 2_c1-
rlabel metal1 -1309 1247 -1309 1247 1 1_c0
rlabel metal1 -1302 1247 -1302 1247 1 1_c0-
rlabel metal1 -1295 1247 -1295 1247 1 1_c1
rlabel metal1 -1288 1247 -1288 1247 1 1_c1-
rlabel metal2 230 1140 230 1140 1 penultimate_bit9
rlabel metal1 347 1252 347 1252 1 last_c0
rlabel metal1 354 1252 354 1252 1 last_c0-
rlabel metal1 361 1252 361 1252 1 last_c1
rlabel metal1 368 1252 368 1252 1 last_c1-
rlabel metal2 232 1017 232 1017 1 penultimate_bit8
rlabel metal2 432 1017 432 1017 1 last_bit8
rlabel metal1 384 1163 384 1163 1 stage_3
rlabel metal1 384 1197 384 1197 1 stage_2
rlabel metal1 392 1224 392 1224 1 stage_1
rlabel metal2 434 74 434 74 1 last_bit0
rlabel metal2 433 198 433 199 1 last_bit1
rlabel metal2 432 321 432 322 1 last_bit2
rlabel metal2 432 446 432 447 1 last_bit3
rlabel metal2 432 569 432 570 1 last_bit4
rlabel metal2 432 693 432 694 1 last_bit5
rlabel metal2 432 817 432 818 1 last_bit6
rlabel metal2 431 941 431 942 1 last_bit7
rlabel space 1041 1364 1041 1364 1 add_latch_control
rlabel metal2 -286 -231 -286 -231 1 64_bit0
rlabel metal2 39 24 39 24 1 16_bit0
rlabel metal2 75 1491 75 1491 1 s1
rlabel metal2 75 1484 75 1484 1 s0
rlabel metal1 -1556 -208 -1556 -208 1 input_latch_control
rlabel metal2 -1579 -1406 -1579 -1406 1 i9
rlabel metal1 -1535 -207 -1535 -207 1 _input_latch_control
rlabel metal1 1688 -212 1688 -212 1 loop_latch_control
rlabel metal1 1652 -214 1652 -214 1 _loop_latch_control
rlabel metal3 598 78 598 78 1 o0
rlabel m3contact 288 1492 288 1492 1 in_latch
rlabel metal2 297 1492 297 1492 1 loop_latch
rlabel metal1 1019 1187 1023 1187 1 sum_bit9
rlabel metal2 1006 1313 1006 1313 1 cout
rlabel metal1 -177 2360 -129 2388 1 t4
rlabel metal1 -1107 2380 -1093 2391 1 t1
<< end >>
