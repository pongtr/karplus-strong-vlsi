magic
tech scmos
timestamp 1509681502
<< ntransistor >>
rect 42 -22 44 -18
rect 42 -38 44 -34
rect 42 -54 44 -50
rect 90 -6 92 -2
rect 90 -30 92 -26
rect 106 -6 108 -2
rect 161 5 165 7
rect 201 5 205 7
rect 122 -6 124 -2
rect 172 -3 176 -1
rect 302 0 312 2
rect 193 -3 197 -1
rect 106 -14 108 -10
rect 114 -14 116 -10
rect 106 -22 108 -18
rect 114 -22 116 -18
rect 106 -30 108 -26
rect 114 -30 116 -26
rect 98 -38 100 -34
rect 90 -46 92 -42
rect 98 -46 100 -42
rect 90 -54 92 -50
rect 98 -54 100 -50
rect 90 -62 92 -58
rect 98 -62 100 -58
rect 82 -70 84 -66
rect 82 -78 84 -74
rect 161 -11 165 -9
rect 371 -3 375 -1
rect 379 -3 383 -1
rect 322 -8 332 -6
rect 537 -3 541 -1
rect 201 -11 205 -9
rect 172 -19 176 -17
rect 379 -11 383 -9
rect 302 -16 312 -14
rect 193 -19 197 -17
rect 161 -27 165 -25
rect 355 -19 359 -17
rect 322 -24 332 -22
rect 201 -27 205 -25
rect 122 -38 124 -34
rect 172 -35 176 -33
rect 427 -27 431 -25
rect 435 -27 439 -25
rect 302 -32 312 -30
rect 193 -35 197 -33
rect 122 -46 124 -42
rect 161 -43 165 -41
rect 114 -54 116 -50
rect 114 -62 116 -58
rect 106 -78 108 -74
rect 347 -35 351 -33
rect 355 -35 359 -33
rect 322 -40 332 -38
rect 201 -43 205 -41
rect 172 -51 176 -49
rect 395 -43 399 -41
rect 302 -48 312 -46
rect 465 -43 469 -41
rect 193 -51 197 -49
rect 161 -59 165 -57
rect 363 -51 367 -49
rect 322 -56 332 -54
rect 201 -59 205 -57
rect 122 -70 124 -66
rect 172 -67 176 -65
rect 379 -59 383 -57
rect 411 -59 415 -57
rect 302 -64 312 -62
rect 481 -59 485 -57
rect 489 -59 493 -57
rect 193 -67 197 -65
rect 122 -78 124 -74
rect 395 -67 399 -65
rect 322 -72 332 -70
rect 42 -117 44 -113
rect 42 -133 44 -129
rect 42 -157 44 -153
rect 58 -157 60 -153
rect 66 -157 68 -153
rect 42 -165 44 -161
rect 50 -165 52 -161
rect 82 -117 84 -113
rect 82 -125 84 -121
rect 82 -133 84 -129
rect 82 -141 84 -137
rect 82 -149 84 -145
rect 74 -165 76 -161
rect 106 -117 108 -113
rect 114 -117 116 -113
rect 106 -125 108 -121
rect 114 -125 116 -121
rect 98 -133 100 -129
rect 98 -141 100 -137
rect 98 -149 100 -145
rect 90 -157 92 -153
rect 90 -165 92 -161
rect 161 -106 165 -104
rect 201 -106 205 -104
rect 172 -114 176 -112
rect 302 -111 312 -109
rect 505 -75 509 -73
rect 193 -114 197 -112
rect 161 -122 165 -120
rect 363 -114 367 -112
rect 322 -119 332 -117
rect 201 -122 205 -120
rect 122 -133 124 -129
rect 172 -130 176 -128
rect 387 -122 391 -120
rect 302 -127 312 -125
rect 513 -122 517 -120
rect 193 -130 197 -128
rect 122 -141 124 -137
rect 161 -138 165 -136
rect 114 -149 116 -145
rect 106 -157 108 -153
rect 106 -165 108 -161
rect 363 -130 367 -128
rect 322 -135 332 -133
rect 201 -138 205 -136
rect 172 -146 176 -144
rect 302 -143 312 -141
rect 521 -138 525 -136
rect 193 -146 197 -144
rect 122 -157 124 -153
rect 419 -146 423 -144
rect 322 -151 332 -149
rect 529 -146 533 -144
rect 201 -154 205 -152
rect 122 -165 124 -161
rect 347 -154 351 -152
rect 302 -159 312 -157
rect 193 -162 197 -160
rect 347 -162 351 -160
rect 363 -162 367 -160
rect 40 -198 42 -185
rect 32 -221 34 -208
rect 56 -198 58 -185
rect 48 -221 50 -208
rect 72 -198 74 -185
rect 64 -221 66 -208
rect 88 -198 90 -185
rect 80 -221 82 -208
rect 104 -198 106 -185
rect 96 -221 98 -208
rect 120 -198 122 -185
rect 360 -195 362 -183
rect 112 -221 114 -208
rect 352 -208 354 -198
rect 376 -195 378 -183
rect 368 -208 370 -198
rect 392 -195 394 -183
rect 384 -208 386 -198
rect 352 -362 354 -350
rect 408 -195 410 -183
rect 400 -208 402 -198
rect 368 -362 370 -350
rect 41 -373 45 -371
rect 57 -373 61 -371
rect 73 -373 77 -371
rect 89 -373 93 -371
rect 105 -373 109 -371
rect 121 -373 125 -371
rect 41 -378 45 -376
rect 57 -378 61 -376
rect 73 -378 77 -376
rect 89 -378 93 -376
rect 105 -378 109 -376
rect 121 -378 125 -376
rect 360 -377 362 -365
rect 424 -195 426 -183
rect 416 -208 418 -198
rect 384 -362 386 -350
rect 376 -377 378 -365
rect 440 -195 442 -183
rect 432 -208 434 -198
rect 400 -362 402 -350
rect 392 -377 394 -365
rect 478 -195 480 -183
rect 470 -208 472 -198
rect 416 -362 418 -350
rect 408 -377 410 -365
rect 494 -195 496 -183
rect 486 -208 488 -198
rect 432 -362 434 -350
rect 424 -377 426 -365
rect 510 -195 512 -183
rect 502 -208 504 -198
rect 470 -362 472 -350
rect 440 -377 442 -365
rect 526 -195 528 -183
rect 518 -208 520 -198
rect 486 -362 488 -350
rect 478 -377 480 -365
rect 542 -195 544 -183
rect 534 -208 536 -198
rect 502 -362 504 -350
rect 494 -377 496 -365
rect 518 -362 520 -350
rect 510 -377 512 -365
rect 534 -362 536 -350
rect 526 -377 528 -365
rect 542 -377 544 -365
<< ptransistor >>
rect 347 21 351 23
rect 355 21 359 23
rect 363 21 367 23
rect 371 21 375 23
rect 379 21 383 23
rect 387 21 391 23
rect 395 21 399 23
rect 403 21 407 23
rect 411 21 415 23
rect 419 21 423 23
rect 427 21 431 23
rect 435 21 439 23
rect 465 21 469 23
rect 473 21 477 23
rect 481 21 485 23
rect 489 21 493 23
rect 497 21 501 23
rect 505 21 509 23
rect 513 21 517 23
rect 521 21 525 23
rect 529 21 533 23
rect 537 21 541 23
rect 10 -6 12 -2
rect 10 -14 12 -10
rect 10 -22 12 -18
rect 10 -30 12 -26
rect 10 -38 12 -34
rect 10 -46 12 -42
rect 10 -54 12 -50
rect 10 -62 12 -58
rect 10 -70 12 -66
rect 10 -78 12 -74
rect 145 5 149 7
rect 217 5 221 7
rect 145 -3 149 -1
rect 270 0 290 2
rect 217 -3 221 -1
rect 145 -11 149 -9
rect 240 -8 260 -6
rect 217 -11 221 -9
rect 145 -19 149 -17
rect 270 -16 290 -14
rect 217 -19 221 -17
rect 145 -27 149 -25
rect 240 -24 260 -22
rect 217 -27 221 -25
rect 145 -35 149 -33
rect 270 -32 290 -30
rect 217 -35 221 -33
rect 145 -43 149 -41
rect 240 -40 260 -38
rect 217 -43 221 -41
rect 145 -51 149 -49
rect 270 -48 290 -46
rect 217 -51 221 -49
rect 145 -59 149 -57
rect 240 -56 260 -54
rect 217 -59 221 -57
rect 145 -67 149 -65
rect 270 -64 290 -62
rect 217 -67 221 -65
rect 240 -72 260 -70
rect 10 -117 12 -113
rect 10 -125 12 -121
rect 10 -133 12 -129
rect 10 -141 12 -137
rect 10 -149 12 -145
rect 10 -157 12 -153
rect 10 -165 12 -161
rect 145 -106 149 -104
rect 217 -106 221 -104
rect 145 -114 149 -112
rect 270 -111 290 -109
rect 217 -114 221 -112
rect 145 -122 149 -120
rect 240 -119 260 -117
rect 217 -122 221 -120
rect 145 -130 149 -128
rect 270 -127 290 -125
rect 217 -130 221 -128
rect 145 -138 149 -136
rect 240 -135 260 -133
rect 217 -138 221 -136
rect 145 -146 149 -144
rect 270 -143 290 -141
rect 217 -146 221 -144
rect 240 -151 260 -149
rect 217 -154 221 -152
rect 270 -159 290 -157
rect 217 -162 221 -160
rect 32 -258 34 -233
rect 48 -258 50 -233
rect 40 -294 42 -268
rect 64 -258 66 -233
rect 56 -294 58 -268
rect 80 -258 82 -233
rect 72 -294 74 -268
rect 96 -258 98 -233
rect 88 -294 90 -268
rect 112 -258 114 -233
rect 104 -294 106 -268
rect 352 -244 354 -220
rect 368 -244 370 -220
rect 120 -294 122 -268
rect 41 -312 45 -310
rect 57 -312 61 -310
rect 73 -312 77 -310
rect 89 -312 93 -310
rect 105 -312 109 -310
rect 121 -312 125 -310
rect 41 -317 45 -315
rect 57 -317 61 -315
rect 73 -317 77 -315
rect 89 -317 93 -315
rect 105 -317 109 -315
rect 121 -317 125 -315
rect 360 -271 362 -247
rect 384 -244 386 -220
rect 360 -312 362 -288
rect 41 -344 45 -342
rect 57 -344 61 -342
rect 73 -344 77 -342
rect 89 -344 93 -342
rect 105 -344 109 -342
rect 352 -338 354 -316
rect 121 -344 125 -342
rect 41 -349 45 -347
rect 57 -349 61 -347
rect 73 -349 77 -347
rect 89 -349 93 -347
rect 105 -349 109 -347
rect 121 -349 125 -347
rect 376 -271 378 -247
rect 400 -244 402 -220
rect 376 -312 378 -288
rect 368 -338 370 -316
rect 392 -271 394 -247
rect 416 -244 418 -220
rect 392 -312 394 -288
rect 384 -338 386 -316
rect 408 -271 410 -247
rect 432 -244 434 -220
rect 408 -312 410 -288
rect 400 -338 402 -316
rect 424 -271 426 -247
rect 470 -244 472 -220
rect 424 -312 426 -288
rect 416 -338 418 -316
rect 440 -271 442 -247
rect 486 -244 488 -220
rect 440 -312 442 -288
rect 432 -338 434 -316
rect 478 -271 480 -247
rect 502 -244 504 -220
rect 478 -312 480 -288
rect 470 -338 472 -316
rect 494 -271 496 -247
rect 518 -244 520 -220
rect 494 -312 496 -288
rect 486 -338 488 -316
rect 510 -271 512 -247
rect 534 -244 536 -220
rect 510 -312 512 -288
rect 502 -338 504 -316
rect 526 -271 528 -247
rect 526 -312 528 -288
rect 518 -338 520 -316
rect 542 -271 544 -247
rect 542 -312 544 -288
rect 534 -338 536 -316
<< ndiffusion >>
rect 37 -18 41 1
rect 37 -22 42 -18
rect 44 -22 45 -18
rect 37 -34 41 -22
rect 37 -38 42 -34
rect 44 -38 45 -34
rect 37 -50 41 -38
rect 37 -54 42 -50
rect 44 -54 45 -50
rect 37 -81 41 -54
rect 53 -81 57 1
rect 69 -81 73 1
rect 85 -2 89 1
rect 85 -6 90 -2
rect 92 -6 93 -2
rect 85 -26 89 -6
rect 85 -30 90 -26
rect 92 -30 93 -26
rect 85 -42 89 -30
rect 101 -2 105 1
rect 101 -6 106 -2
rect 108 -6 109 -2
rect 101 -10 105 -6
rect 117 -2 121 1
rect 161 7 165 8
rect 161 3 165 5
rect 201 7 205 8
rect 201 3 205 5
rect 161 0 176 3
rect 172 -1 176 0
rect 117 -6 122 -2
rect 124 -6 125 -2
rect 193 0 205 3
rect 193 -1 197 0
rect 302 2 312 3
rect 117 -10 121 -6
rect 101 -14 106 -10
rect 108 -14 109 -10
rect 113 -14 114 -10
rect 116 -14 121 -10
rect 101 -18 105 -14
rect 117 -18 121 -14
rect 101 -22 106 -18
rect 108 -22 109 -18
rect 113 -22 114 -18
rect 116 -22 121 -18
rect 101 -26 105 -22
rect 117 -26 121 -22
rect 101 -30 106 -26
rect 108 -30 109 -26
rect 113 -30 114 -26
rect 116 -30 121 -26
rect 101 -34 105 -30
rect 97 -38 98 -34
rect 100 -38 105 -34
rect 101 -42 105 -38
rect 85 -46 90 -42
rect 92 -46 93 -42
rect 97 -46 98 -42
rect 100 -46 105 -42
rect 85 -50 89 -46
rect 101 -50 105 -46
rect 85 -54 90 -50
rect 92 -54 93 -50
rect 97 -54 98 -50
rect 100 -54 105 -50
rect 85 -58 89 -54
rect 101 -58 105 -54
rect 85 -62 90 -58
rect 92 -62 93 -58
rect 97 -62 98 -58
rect 100 -62 105 -58
rect 85 -66 89 -62
rect 81 -70 82 -66
rect 84 -70 89 -66
rect 85 -74 89 -70
rect 81 -78 82 -74
rect 84 -78 89 -74
rect 85 -81 89 -78
rect 101 -74 105 -62
rect 117 -34 121 -30
rect 172 -4 176 -3
rect 193 -4 197 -3
rect 172 -7 175 -4
rect 161 -9 165 -8
rect 161 -13 165 -11
rect 201 -9 205 -8
rect 302 -1 312 0
rect 371 -1 375 0
rect 379 -1 383 0
rect 537 -1 541 0
rect 314 -5 315 -1
rect 319 -5 320 -1
rect 330 -5 332 -1
rect 371 -4 375 -3
rect 379 -4 383 -3
rect 322 -6 332 -5
rect 343 -8 444 -4
rect 537 -4 541 -3
rect 461 -8 546 -4
rect 322 -9 332 -8
rect 379 -9 383 -8
rect 201 -13 205 -11
rect 161 -16 176 -13
rect 172 -17 176 -16
rect 193 -16 205 -13
rect 193 -17 197 -16
rect 379 -12 383 -11
rect 302 -14 312 -13
rect 172 -20 176 -19
rect 193 -20 197 -19
rect 172 -23 175 -20
rect 161 -25 165 -24
rect 161 -29 165 -27
rect 201 -25 205 -24
rect 302 -17 312 -16
rect 355 -17 359 -16
rect 314 -21 315 -17
rect 319 -21 320 -17
rect 330 -21 332 -17
rect 355 -20 359 -19
rect 322 -22 332 -21
rect 343 -24 444 -20
rect 461 -24 546 -20
rect 322 -25 332 -24
rect 427 -25 431 -24
rect 435 -25 439 -24
rect 201 -29 205 -27
rect 161 -32 176 -29
rect 172 -33 176 -32
rect 117 -38 122 -34
rect 124 -38 125 -34
rect 193 -32 205 -29
rect 193 -33 197 -32
rect 427 -28 431 -27
rect 302 -30 312 -29
rect 117 -42 121 -38
rect 117 -46 122 -42
rect 124 -46 125 -42
rect 172 -36 176 -35
rect 193 -36 197 -35
rect 172 -39 175 -36
rect 161 -41 165 -40
rect 117 -50 121 -46
rect 113 -54 114 -50
rect 116 -54 121 -50
rect 117 -58 121 -54
rect 113 -62 114 -58
rect 116 -62 121 -58
rect 101 -78 106 -74
rect 108 -78 109 -74
rect 101 -81 105 -78
rect 117 -66 121 -62
rect 161 -45 165 -43
rect 201 -41 205 -40
rect 302 -33 312 -32
rect 347 -33 351 -32
rect 435 -28 439 -27
rect 355 -33 359 -32
rect 314 -37 315 -33
rect 319 -37 320 -33
rect 330 -37 332 -33
rect 347 -36 351 -35
rect 355 -36 359 -35
rect 322 -38 332 -37
rect 343 -40 444 -36
rect 461 -40 546 -36
rect 322 -41 332 -40
rect 395 -41 399 -40
rect 465 -41 469 -40
rect 201 -45 205 -43
rect 161 -48 176 -45
rect 172 -49 176 -48
rect 193 -48 205 -45
rect 193 -49 197 -48
rect 395 -44 399 -43
rect 302 -46 312 -45
rect 465 -44 469 -43
rect 172 -52 176 -51
rect 193 -52 197 -51
rect 172 -55 175 -52
rect 161 -57 165 -56
rect 161 -61 165 -59
rect 201 -57 205 -56
rect 302 -49 312 -48
rect 363 -49 367 -48
rect 314 -53 315 -49
rect 319 -53 320 -49
rect 330 -53 332 -49
rect 363 -52 367 -51
rect 322 -54 332 -53
rect 343 -56 444 -52
rect 461 -56 546 -52
rect 322 -57 332 -56
rect 379 -57 383 -56
rect 411 -57 415 -56
rect 481 -57 485 -56
rect 489 -57 493 -56
rect 201 -61 205 -59
rect 161 -64 176 -61
rect 172 -65 176 -64
rect 117 -70 122 -66
rect 124 -70 125 -66
rect 193 -64 205 -61
rect 193 -65 197 -64
rect 379 -60 383 -59
rect 411 -60 415 -59
rect 302 -62 312 -61
rect 481 -60 485 -59
rect 489 -60 493 -59
rect 117 -74 121 -70
rect 117 -78 122 -74
rect 124 -78 125 -74
rect 172 -68 176 -67
rect 193 -68 197 -67
rect 172 -71 175 -68
rect 302 -65 312 -64
rect 395 -65 399 -64
rect 314 -69 315 -65
rect 319 -69 320 -65
rect 330 -69 332 -65
rect 395 -68 399 -67
rect 322 -70 332 -69
rect 343 -72 444 -68
rect 461 -72 546 -68
rect 322 -73 332 -72
rect 505 -73 509 -72
rect 117 -81 121 -78
rect 37 -113 41 -110
rect 37 -117 42 -113
rect 44 -117 45 -113
rect 37 -129 41 -117
rect 37 -133 42 -129
rect 44 -133 45 -129
rect 37 -153 41 -133
rect 37 -157 42 -153
rect 44 -157 45 -153
rect 37 -161 41 -157
rect 53 -153 57 -110
rect 69 -153 73 -110
rect 53 -157 58 -153
rect 60 -157 61 -153
rect 65 -157 66 -153
rect 68 -157 73 -153
rect 53 -161 57 -157
rect 37 -165 42 -161
rect 44 -165 45 -161
rect 49 -165 50 -161
rect 52 -165 57 -161
rect 37 -168 41 -165
rect 53 -168 57 -165
rect 69 -161 73 -157
rect 85 -113 89 -110
rect 81 -117 82 -113
rect 84 -117 89 -113
rect 85 -121 89 -117
rect 81 -125 82 -121
rect 84 -125 89 -121
rect 85 -129 89 -125
rect 81 -133 82 -129
rect 84 -133 89 -129
rect 85 -137 89 -133
rect 81 -141 82 -137
rect 84 -141 89 -137
rect 85 -145 89 -141
rect 81 -149 82 -145
rect 84 -149 89 -145
rect 69 -165 74 -161
rect 76 -165 77 -161
rect 69 -168 73 -165
rect 85 -153 89 -149
rect 101 -113 105 -110
rect 117 -113 121 -110
rect 101 -117 106 -113
rect 108 -117 109 -113
rect 113 -117 114 -113
rect 116 -117 121 -113
rect 101 -121 105 -117
rect 117 -121 121 -117
rect 101 -125 106 -121
rect 108 -125 109 -121
rect 113 -125 114 -121
rect 116 -125 121 -121
rect 101 -129 105 -125
rect 97 -133 98 -129
rect 100 -133 105 -129
rect 101 -137 105 -133
rect 97 -141 98 -137
rect 100 -141 105 -137
rect 101 -145 105 -141
rect 97 -149 98 -145
rect 100 -149 105 -145
rect 85 -157 90 -153
rect 92 -157 93 -153
rect 85 -161 89 -157
rect 85 -165 90 -161
rect 92 -165 93 -161
rect 85 -168 89 -165
rect 101 -153 105 -149
rect 117 -129 121 -125
rect 161 -104 165 -103
rect 161 -108 165 -106
rect 201 -104 205 -103
rect 201 -108 205 -106
rect 161 -111 176 -108
rect 172 -112 176 -111
rect 193 -111 205 -108
rect 193 -112 197 -111
rect 302 -109 312 -108
rect 505 -76 509 -75
rect 172 -115 176 -114
rect 193 -115 197 -114
rect 172 -118 175 -115
rect 161 -120 165 -119
rect 161 -124 165 -122
rect 201 -120 205 -119
rect 302 -112 312 -111
rect 363 -112 367 -111
rect 314 -116 315 -112
rect 319 -116 320 -112
rect 330 -116 332 -112
rect 363 -115 367 -114
rect 322 -117 332 -116
rect 343 -119 444 -115
rect 461 -119 546 -115
rect 322 -120 332 -119
rect 387 -120 391 -119
rect 513 -120 517 -119
rect 201 -124 205 -122
rect 161 -127 176 -124
rect 172 -128 176 -127
rect 117 -133 122 -129
rect 124 -133 125 -129
rect 193 -127 205 -124
rect 193 -128 197 -127
rect 387 -123 391 -122
rect 302 -125 312 -124
rect 513 -123 517 -122
rect 117 -137 121 -133
rect 117 -141 122 -137
rect 124 -141 125 -137
rect 172 -131 176 -130
rect 193 -131 197 -130
rect 172 -134 175 -131
rect 161 -136 165 -135
rect 117 -145 121 -141
rect 113 -149 114 -145
rect 116 -149 121 -145
rect 101 -157 106 -153
rect 108 -157 109 -153
rect 101 -161 105 -157
rect 101 -165 106 -161
rect 108 -165 109 -161
rect 101 -168 105 -165
rect 117 -153 121 -149
rect 161 -140 165 -138
rect 201 -136 205 -135
rect 302 -128 312 -127
rect 363 -128 367 -127
rect 314 -132 315 -128
rect 319 -132 320 -128
rect 330 -132 332 -128
rect 363 -131 367 -130
rect 322 -133 332 -132
rect 343 -135 444 -131
rect 461 -135 546 -131
rect 322 -136 332 -135
rect 521 -136 525 -135
rect 201 -140 205 -138
rect 161 -143 176 -140
rect 172 -144 176 -143
rect 193 -143 205 -140
rect 193 -144 197 -143
rect 302 -141 312 -140
rect 521 -139 525 -138
rect 117 -157 122 -153
rect 124 -157 125 -153
rect 172 -147 176 -146
rect 193 -147 197 -146
rect 172 -150 175 -147
rect 201 -152 205 -151
rect 302 -144 312 -143
rect 419 -144 423 -143
rect 529 -144 533 -143
rect 314 -148 315 -144
rect 319 -148 320 -144
rect 330 -148 332 -144
rect 419 -147 423 -146
rect 322 -149 332 -148
rect 343 -151 444 -147
rect 529 -147 533 -146
rect 461 -151 546 -147
rect 322 -152 332 -151
rect 347 -152 351 -151
rect 201 -156 205 -154
rect 117 -161 121 -157
rect 117 -165 122 -161
rect 124 -165 125 -161
rect 193 -159 205 -156
rect 193 -160 197 -159
rect 347 -155 351 -154
rect 302 -157 312 -156
rect 193 -163 197 -162
rect 117 -168 121 -165
rect 302 -160 312 -159
rect 347 -160 351 -159
rect 363 -160 367 -159
rect 314 -164 315 -160
rect 347 -163 351 -162
rect 363 -163 367 -162
rect 343 -167 444 -163
rect 461 -167 546 -163
rect 363 -181 367 -180
rect 37 -187 40 -185
rect 39 -198 40 -187
rect 42 -198 43 -185
rect 53 -187 56 -185
rect 35 -201 39 -200
rect 35 -206 39 -205
rect 31 -221 32 -208
rect 34 -221 35 -208
rect 55 -198 56 -187
rect 58 -198 59 -185
rect 69 -187 72 -185
rect 51 -201 55 -200
rect 51 -206 55 -205
rect 47 -221 48 -208
rect 50 -221 51 -208
rect 71 -198 72 -187
rect 74 -198 75 -185
rect 85 -187 88 -185
rect 67 -201 71 -200
rect 67 -206 71 -205
rect 63 -221 64 -208
rect 66 -221 67 -208
rect 87 -198 88 -187
rect 90 -198 91 -185
rect 101 -187 104 -185
rect 83 -201 87 -200
rect 83 -206 87 -205
rect 79 -221 80 -208
rect 82 -221 83 -208
rect 103 -198 104 -187
rect 106 -198 107 -185
rect 117 -187 120 -185
rect 99 -201 103 -200
rect 99 -206 103 -205
rect 95 -221 96 -208
rect 98 -221 99 -208
rect 119 -198 120 -187
rect 122 -198 123 -185
rect 356 -195 360 -183
rect 362 -190 363 -183
rect 379 -181 383 -180
rect 362 -195 366 -190
rect 356 -198 359 -195
rect 115 -201 119 -200
rect 115 -206 119 -205
rect 111 -221 112 -208
rect 114 -221 115 -208
rect 348 -200 352 -198
rect 351 -208 352 -200
rect 354 -208 359 -198
rect 372 -195 376 -183
rect 378 -190 379 -183
rect 395 -181 399 -180
rect 378 -195 382 -190
rect 372 -198 375 -195
rect 364 -200 368 -198
rect 367 -208 368 -200
rect 370 -208 375 -198
rect 388 -195 392 -183
rect 394 -190 395 -183
rect 411 -181 415 -180
rect 394 -195 398 -190
rect 388 -198 391 -195
rect 380 -200 384 -198
rect 383 -208 384 -200
rect 386 -208 391 -198
rect 351 -360 352 -350
rect 348 -362 352 -360
rect 354 -362 359 -350
rect 47 -370 48 -366
rect 41 -371 45 -370
rect 63 -370 64 -366
rect 57 -371 61 -370
rect 79 -370 80 -366
rect 73 -371 77 -370
rect 95 -370 96 -366
rect 89 -371 93 -370
rect 111 -370 112 -366
rect 105 -371 109 -370
rect 127 -370 128 -366
rect 356 -365 359 -362
rect 404 -195 408 -183
rect 410 -190 411 -183
rect 427 -181 431 -180
rect 410 -195 414 -190
rect 404 -198 407 -195
rect 396 -200 400 -198
rect 399 -208 400 -200
rect 402 -208 407 -198
rect 367 -360 368 -350
rect 364 -362 368 -360
rect 370 -362 375 -350
rect 121 -371 125 -370
rect 41 -376 45 -373
rect 57 -376 61 -373
rect 73 -376 77 -373
rect 89 -376 93 -373
rect 105 -376 109 -373
rect 121 -376 125 -373
rect 41 -379 45 -378
rect 41 -382 42 -379
rect 57 -379 61 -378
rect 57 -382 58 -379
rect 73 -379 77 -378
rect 73 -382 74 -379
rect 89 -379 93 -378
rect 89 -382 90 -379
rect 105 -379 109 -378
rect 105 -382 106 -379
rect 356 -377 360 -365
rect 362 -370 366 -365
rect 372 -365 375 -362
rect 420 -195 424 -183
rect 426 -190 427 -183
rect 443 -181 447 -180
rect 426 -195 430 -190
rect 420 -198 423 -195
rect 412 -200 416 -198
rect 415 -208 416 -200
rect 418 -208 423 -198
rect 383 -360 384 -350
rect 380 -362 384 -360
rect 386 -362 391 -350
rect 362 -377 363 -370
rect 121 -379 125 -378
rect 372 -377 376 -365
rect 378 -370 382 -365
rect 388 -365 391 -362
rect 436 -195 440 -183
rect 442 -190 443 -183
rect 481 -181 485 -180
rect 442 -195 446 -190
rect 436 -198 439 -195
rect 428 -200 432 -198
rect 431 -208 432 -200
rect 434 -208 439 -198
rect 399 -360 400 -350
rect 396 -362 400 -360
rect 402 -362 407 -350
rect 378 -377 379 -370
rect 388 -377 392 -365
rect 394 -370 398 -365
rect 404 -365 407 -362
rect 474 -195 478 -183
rect 480 -190 481 -183
rect 497 -181 501 -180
rect 480 -195 484 -190
rect 474 -198 477 -195
rect 466 -200 470 -198
rect 469 -208 470 -200
rect 472 -208 477 -198
rect 415 -360 416 -350
rect 412 -362 416 -360
rect 418 -362 423 -350
rect 394 -377 395 -370
rect 404 -377 408 -365
rect 410 -370 414 -365
rect 420 -365 423 -362
rect 490 -195 494 -183
rect 496 -190 497 -183
rect 513 -181 517 -180
rect 496 -195 500 -190
rect 490 -198 493 -195
rect 482 -200 486 -198
rect 485 -208 486 -200
rect 488 -208 493 -198
rect 431 -360 432 -350
rect 428 -362 432 -360
rect 434 -362 439 -350
rect 410 -377 411 -370
rect 420 -377 424 -365
rect 426 -370 430 -365
rect 436 -365 439 -362
rect 506 -195 510 -183
rect 512 -190 513 -183
rect 529 -181 533 -180
rect 512 -195 516 -190
rect 506 -198 509 -195
rect 498 -200 502 -198
rect 501 -208 502 -200
rect 504 -208 509 -198
rect 469 -360 470 -350
rect 466 -362 470 -360
rect 472 -362 477 -350
rect 426 -377 427 -370
rect 436 -377 440 -365
rect 442 -370 446 -365
rect 474 -365 477 -362
rect 522 -195 526 -183
rect 528 -190 529 -183
rect 545 -181 549 -180
rect 528 -195 532 -190
rect 522 -198 525 -195
rect 514 -200 518 -198
rect 517 -208 518 -200
rect 520 -208 525 -198
rect 485 -360 486 -350
rect 482 -362 486 -360
rect 488 -362 493 -350
rect 442 -377 443 -370
rect 474 -377 478 -365
rect 480 -370 484 -365
rect 490 -365 493 -362
rect 538 -195 542 -183
rect 544 -190 545 -183
rect 544 -195 548 -190
rect 538 -198 541 -195
rect 530 -200 534 -198
rect 533 -208 534 -200
rect 536 -208 541 -198
rect 501 -360 502 -350
rect 498 -362 502 -360
rect 504 -362 509 -350
rect 480 -377 481 -370
rect 490 -377 494 -365
rect 496 -370 500 -365
rect 506 -365 509 -362
rect 517 -360 518 -350
rect 514 -362 518 -360
rect 520 -362 525 -350
rect 496 -377 497 -370
rect 506 -377 510 -365
rect 512 -370 516 -365
rect 522 -365 525 -362
rect 533 -360 534 -350
rect 530 -362 534 -360
rect 536 -362 541 -350
rect 512 -377 513 -370
rect 522 -377 526 -365
rect 528 -370 532 -365
rect 538 -365 541 -362
rect 528 -377 529 -370
rect 538 -377 542 -365
rect 544 -370 548 -365
rect 544 -377 545 -370
rect 121 -382 122 -379
rect 363 -380 367 -379
rect 379 -380 383 -379
rect 395 -380 399 -379
rect 411 -380 415 -379
rect 427 -380 431 -379
rect 443 -380 447 -379
rect 481 -380 485 -379
rect 497 -380 501 -379
rect 513 -380 517 -379
rect 529 -380 533 -379
rect 545 -380 549 -379
<< pdiffusion >>
rect 345 28 543 29
rect 347 23 351 24
rect 355 23 359 24
rect 363 23 367 24
rect 371 23 375 24
rect 379 23 383 24
rect 387 23 391 24
rect 395 23 399 24
rect 403 23 407 24
rect 411 23 415 24
rect 419 23 423 24
rect 427 23 431 24
rect 435 23 439 24
rect 465 23 469 24
rect 473 23 477 24
rect 481 23 485 24
rect 489 23 493 24
rect 497 23 501 24
rect 505 23 509 24
rect 513 23 517 24
rect 521 23 525 24
rect 529 23 533 24
rect 537 23 541 24
rect 347 20 351 21
rect 355 20 359 21
rect 363 20 367 21
rect 371 20 375 21
rect 379 20 383 21
rect 387 20 391 21
rect 395 20 399 21
rect 403 20 407 21
rect 411 20 415 21
rect 419 20 423 21
rect 427 20 431 21
rect 435 20 439 21
rect 465 20 469 21
rect 473 20 477 21
rect 481 20 485 21
rect 489 20 493 21
rect 497 20 501 21
rect 505 20 509 21
rect 513 20 517 21
rect 521 20 525 21
rect 529 20 533 21
rect 537 20 541 21
rect 142 8 143 12
rect 4 -80 5 0
rect 9 -6 10 -2
rect 12 -6 13 -2
rect 9 -14 10 -10
rect 12 -14 13 -10
rect 9 -22 10 -18
rect 12 -22 13 -18
rect 9 -30 10 -26
rect 12 -30 13 -26
rect 9 -38 10 -34
rect 12 -38 13 -34
rect 9 -46 10 -42
rect 12 -46 13 -42
rect 9 -54 10 -50
rect 12 -54 13 -50
rect 9 -62 10 -58
rect 12 -62 13 -58
rect 9 -70 10 -66
rect 12 -70 13 -66
rect 9 -78 10 -74
rect 12 -78 13 -74
rect 145 7 149 8
rect 145 4 149 5
rect 223 8 224 12
rect 217 7 221 8
rect 145 -1 149 0
rect 217 4 221 5
rect 270 3 275 7
rect 217 -1 221 0
rect 270 2 290 3
rect 270 -1 290 0
rect 145 -4 149 -3
rect 217 -4 221 -3
rect 142 -8 143 -4
rect 145 -9 149 -8
rect 145 -12 149 -11
rect 223 -8 224 -4
rect 240 -5 242 -1
rect 262 -5 263 -1
rect 267 -5 268 -1
rect 217 -9 221 -8
rect 240 -6 260 -5
rect 240 -9 260 -8
rect 145 -17 149 -16
rect 217 -12 221 -11
rect 240 -13 242 -9
rect 270 -13 275 -9
rect 217 -17 221 -16
rect 270 -14 290 -13
rect 270 -17 290 -16
rect 145 -20 149 -19
rect 217 -20 221 -19
rect 142 -24 143 -20
rect 145 -25 149 -24
rect 145 -28 149 -27
rect 223 -24 224 -20
rect 240 -21 242 -17
rect 262 -21 263 -17
rect 267 -21 268 -17
rect 217 -25 221 -24
rect 240 -22 260 -21
rect 240 -25 260 -24
rect 145 -33 149 -32
rect 217 -28 221 -27
rect 240 -29 242 -25
rect 270 -29 275 -25
rect 217 -33 221 -32
rect 270 -30 290 -29
rect 270 -33 290 -32
rect 145 -36 149 -35
rect 217 -36 221 -35
rect 142 -40 143 -36
rect 145 -41 149 -40
rect 145 -44 149 -43
rect 223 -40 224 -36
rect 240 -37 242 -33
rect 262 -37 263 -33
rect 267 -37 268 -33
rect 217 -41 221 -40
rect 240 -38 260 -37
rect 240 -41 260 -40
rect 145 -49 149 -48
rect 217 -44 221 -43
rect 240 -45 242 -41
rect 270 -45 275 -41
rect 217 -49 221 -48
rect 270 -46 290 -45
rect 270 -49 290 -48
rect 145 -52 149 -51
rect 217 -52 221 -51
rect 142 -56 143 -52
rect 145 -57 149 -56
rect 145 -60 149 -59
rect 223 -56 224 -52
rect 240 -53 242 -49
rect 262 -53 263 -49
rect 267 -53 268 -49
rect 217 -57 221 -56
rect 240 -54 260 -53
rect 240 -57 260 -56
rect 145 -65 149 -64
rect 217 -60 221 -59
rect 240 -61 242 -57
rect 270 -61 275 -57
rect 217 -65 221 -64
rect 270 -62 290 -61
rect 270 -65 290 -64
rect 145 -68 149 -67
rect 142 -72 143 -68
rect 217 -68 221 -67
rect 223 -72 224 -68
rect 240 -69 242 -65
rect 262 -69 263 -65
rect 267 -69 268 -65
rect 240 -70 260 -69
rect 240 -73 260 -72
rect 240 -77 242 -73
rect 4 -167 5 -111
rect 9 -117 10 -113
rect 12 -117 13 -113
rect 9 -125 10 -121
rect 12 -125 13 -121
rect 9 -133 10 -129
rect 12 -133 13 -129
rect 9 -141 10 -137
rect 12 -141 13 -137
rect 9 -149 10 -145
rect 12 -149 13 -145
rect 9 -157 10 -153
rect 12 -157 13 -153
rect 9 -165 10 -161
rect 12 -165 13 -161
rect 142 -103 143 -99
rect 145 -104 149 -103
rect 145 -107 149 -106
rect 223 -103 224 -99
rect 217 -104 221 -103
rect 145 -112 149 -111
rect 217 -107 221 -106
rect 270 -108 275 -104
rect 217 -112 221 -111
rect 270 -109 290 -108
rect 270 -112 290 -111
rect 145 -115 149 -114
rect 217 -115 221 -114
rect 142 -119 143 -115
rect 145 -120 149 -119
rect 145 -123 149 -122
rect 223 -119 224 -115
rect 240 -116 242 -112
rect 262 -116 263 -112
rect 267 -116 268 -112
rect 217 -120 221 -119
rect 240 -117 260 -116
rect 240 -120 260 -119
rect 145 -128 149 -127
rect 217 -123 221 -122
rect 240 -124 242 -120
rect 270 -124 275 -120
rect 217 -128 221 -127
rect 270 -125 290 -124
rect 270 -128 290 -127
rect 145 -131 149 -130
rect 217 -131 221 -130
rect 142 -135 143 -131
rect 145 -136 149 -135
rect 145 -139 149 -138
rect 223 -135 224 -131
rect 240 -132 242 -128
rect 262 -132 263 -128
rect 267 -132 268 -128
rect 217 -136 221 -135
rect 240 -133 260 -132
rect 240 -136 260 -135
rect 145 -144 149 -143
rect 217 -139 221 -138
rect 240 -140 242 -136
rect 270 -140 275 -136
rect 217 -144 221 -143
rect 270 -141 290 -140
rect 270 -144 290 -143
rect 145 -147 149 -146
rect 142 -151 143 -147
rect 217 -147 221 -146
rect 223 -151 224 -147
rect 240 -148 242 -144
rect 262 -148 263 -144
rect 267 -148 268 -144
rect 217 -152 221 -151
rect 240 -149 260 -148
rect 240 -152 260 -151
rect 217 -155 221 -154
rect 240 -156 242 -152
rect 270 -156 275 -152
rect 217 -160 221 -159
rect 270 -157 290 -156
rect 270 -160 290 -159
rect 217 -163 221 -162
rect 223 -167 224 -163
rect 267 -164 268 -160
rect 31 -251 32 -233
rect 29 -258 32 -251
rect 34 -258 35 -233
rect 35 -261 39 -260
rect 35 -266 39 -265
rect 47 -251 48 -233
rect 45 -258 48 -251
rect 50 -258 51 -233
rect 39 -292 40 -268
rect 35 -294 40 -292
rect 42 -285 43 -268
rect 42 -294 45 -285
rect 51 -261 55 -260
rect 51 -266 55 -265
rect 63 -251 64 -233
rect 61 -258 64 -251
rect 66 -258 67 -233
rect 55 -292 56 -268
rect 51 -294 56 -292
rect 58 -285 59 -268
rect 58 -294 61 -285
rect 67 -261 71 -260
rect 67 -266 71 -265
rect 79 -251 80 -233
rect 77 -258 80 -251
rect 82 -258 83 -233
rect 71 -292 72 -268
rect 67 -294 72 -292
rect 74 -285 75 -268
rect 74 -294 77 -285
rect 83 -261 87 -260
rect 83 -266 87 -265
rect 95 -251 96 -233
rect 93 -258 96 -251
rect 98 -258 99 -233
rect 87 -292 88 -268
rect 83 -294 88 -292
rect 90 -285 91 -268
rect 90 -294 93 -285
rect 99 -261 103 -260
rect 99 -266 103 -265
rect 111 -251 112 -233
rect 109 -258 112 -251
rect 114 -258 115 -233
rect 103 -292 104 -268
rect 99 -294 104 -292
rect 106 -285 107 -268
rect 106 -294 109 -285
rect 115 -261 119 -260
rect 115 -266 119 -265
rect 351 -242 352 -220
rect 348 -244 352 -242
rect 354 -244 359 -220
rect 356 -247 359 -244
rect 367 -242 368 -220
rect 364 -244 368 -242
rect 370 -244 375 -220
rect 119 -292 120 -268
rect 115 -294 120 -292
rect 122 -285 123 -268
rect 122 -294 125 -285
rect 41 -309 42 -307
rect 41 -310 45 -309
rect 57 -309 58 -307
rect 57 -310 61 -309
rect 73 -309 74 -307
rect 73 -310 77 -309
rect 89 -309 90 -307
rect 89 -310 93 -309
rect 105 -309 106 -307
rect 105 -310 109 -309
rect 121 -309 122 -307
rect 121 -310 125 -309
rect 41 -315 45 -312
rect 57 -315 61 -312
rect 73 -315 77 -312
rect 89 -315 93 -312
rect 105 -315 109 -312
rect 121 -315 125 -312
rect 356 -271 360 -247
rect 362 -252 366 -247
rect 372 -247 375 -244
rect 383 -242 384 -220
rect 380 -244 384 -242
rect 386 -244 391 -220
rect 362 -271 363 -252
rect 363 -274 367 -273
rect 356 -312 360 -288
rect 362 -312 363 -288
rect 356 -316 359 -312
rect 41 -318 45 -317
rect 47 -322 48 -318
rect 57 -318 61 -317
rect 63 -322 64 -318
rect 73 -318 77 -317
rect 79 -322 80 -318
rect 89 -318 93 -317
rect 95 -322 96 -318
rect 105 -318 109 -317
rect 111 -322 112 -318
rect 121 -318 125 -317
rect 127 -322 128 -318
rect 41 -341 42 -339
rect 41 -342 45 -341
rect 57 -341 58 -339
rect 57 -342 61 -341
rect 73 -341 74 -339
rect 73 -342 77 -341
rect 89 -341 90 -339
rect 89 -342 93 -341
rect 105 -341 106 -339
rect 105 -342 109 -341
rect 121 -341 122 -339
rect 351 -338 352 -316
rect 354 -338 359 -316
rect 121 -342 125 -341
rect 41 -347 45 -344
rect 57 -347 61 -344
rect 73 -347 77 -344
rect 89 -347 93 -344
rect 105 -347 109 -344
rect 121 -347 125 -344
rect 41 -350 45 -349
rect 47 -354 48 -350
rect 57 -350 61 -349
rect 63 -354 64 -350
rect 73 -350 77 -349
rect 79 -354 80 -350
rect 89 -350 93 -349
rect 95 -354 96 -350
rect 105 -350 109 -349
rect 111 -354 112 -350
rect 121 -350 125 -349
rect 127 -354 128 -350
rect 372 -271 376 -247
rect 378 -252 382 -247
rect 388 -247 391 -244
rect 399 -242 400 -220
rect 396 -244 400 -242
rect 402 -244 407 -220
rect 378 -271 379 -252
rect 379 -274 383 -273
rect 372 -312 376 -288
rect 378 -312 379 -288
rect 372 -316 375 -312
rect 367 -338 368 -316
rect 370 -338 375 -316
rect 388 -271 392 -247
rect 394 -252 398 -247
rect 404 -247 407 -244
rect 415 -242 416 -220
rect 412 -244 416 -242
rect 418 -244 423 -220
rect 394 -271 395 -252
rect 395 -274 399 -273
rect 388 -312 392 -288
rect 394 -312 395 -288
rect 388 -316 391 -312
rect 383 -338 384 -316
rect 386 -338 391 -316
rect 404 -271 408 -247
rect 410 -252 414 -247
rect 420 -247 423 -244
rect 431 -242 432 -220
rect 428 -244 432 -242
rect 434 -244 439 -220
rect 410 -271 411 -252
rect 411 -274 415 -273
rect 404 -312 408 -288
rect 410 -312 411 -288
rect 404 -316 407 -312
rect 399 -338 400 -316
rect 402 -338 407 -316
rect 420 -271 424 -247
rect 426 -252 430 -247
rect 436 -247 439 -244
rect 469 -242 470 -220
rect 466 -244 470 -242
rect 472 -244 477 -220
rect 426 -271 427 -252
rect 427 -274 431 -273
rect 420 -312 424 -288
rect 426 -312 427 -288
rect 420 -316 423 -312
rect 415 -338 416 -316
rect 418 -338 423 -316
rect 436 -271 440 -247
rect 442 -252 446 -247
rect 474 -247 477 -244
rect 485 -242 486 -220
rect 482 -244 486 -242
rect 488 -244 493 -220
rect 442 -271 443 -252
rect 443 -274 447 -273
rect 436 -312 440 -288
rect 442 -312 443 -288
rect 436 -316 439 -312
rect 431 -338 432 -316
rect 434 -338 439 -316
rect 474 -271 478 -247
rect 480 -252 484 -247
rect 490 -247 493 -244
rect 501 -242 502 -220
rect 498 -244 502 -242
rect 504 -244 509 -220
rect 480 -271 481 -252
rect 481 -274 485 -273
rect 474 -312 478 -288
rect 480 -312 481 -288
rect 474 -316 477 -312
rect 469 -338 470 -316
rect 472 -338 477 -316
rect 490 -271 494 -247
rect 496 -252 500 -247
rect 506 -247 509 -244
rect 517 -242 518 -220
rect 514 -244 518 -242
rect 520 -244 525 -220
rect 496 -271 497 -252
rect 497 -274 501 -273
rect 490 -312 494 -288
rect 496 -312 497 -288
rect 490 -316 493 -312
rect 485 -338 486 -316
rect 488 -338 493 -316
rect 506 -271 510 -247
rect 512 -252 516 -247
rect 522 -247 525 -244
rect 533 -242 534 -220
rect 530 -244 534 -242
rect 536 -244 541 -220
rect 512 -271 513 -252
rect 513 -274 517 -273
rect 506 -312 510 -288
rect 512 -312 513 -288
rect 506 -316 509 -312
rect 501 -338 502 -316
rect 504 -338 509 -316
rect 522 -271 526 -247
rect 528 -252 532 -247
rect 538 -247 541 -244
rect 528 -271 529 -252
rect 529 -274 533 -273
rect 522 -312 526 -288
rect 528 -312 529 -288
rect 522 -316 525 -312
rect 517 -338 518 -316
rect 520 -338 525 -316
rect 538 -271 542 -247
rect 544 -252 548 -247
rect 544 -271 545 -252
rect 545 -274 549 -273
rect 538 -312 542 -288
rect 544 -312 545 -288
rect 538 -316 541 -312
rect 533 -338 534 -316
rect 536 -338 541 -316
<< ndcontact >>
rect 37 1 41 5
rect 45 -22 49 -18
rect 45 -38 49 -34
rect 45 -54 49 -50
rect 37 -85 41 -81
rect 53 1 57 5
rect 53 -85 57 -81
rect 69 1 73 5
rect 69 -85 73 -81
rect 85 1 89 5
rect 93 -6 97 -2
rect 93 -30 97 -26
rect 101 1 105 5
rect 109 -6 113 -2
rect 117 1 121 5
rect 161 8 165 12
rect 201 8 205 12
rect 125 -6 129 -2
rect 302 3 312 7
rect 371 0 375 4
rect 109 -14 113 -10
rect 109 -22 113 -18
rect 109 -30 113 -26
rect 93 -38 97 -34
rect 93 -46 97 -42
rect 93 -54 97 -50
rect 93 -62 97 -58
rect 77 -70 81 -66
rect 77 -78 81 -74
rect 85 -85 89 -81
rect 161 -8 165 -4
rect 175 -8 179 -4
rect 193 -8 197 -4
rect 201 -8 205 -4
rect 379 0 383 4
rect 537 0 541 4
rect 302 -5 314 -1
rect 320 -5 330 -1
rect 444 -8 448 -4
rect 546 -8 550 -4
rect 302 -13 312 -9
rect 322 -13 332 -9
rect 355 -16 359 -12
rect 379 -16 383 -12
rect 161 -24 165 -20
rect 175 -24 179 -20
rect 193 -24 197 -20
rect 201 -24 205 -20
rect 302 -21 314 -17
rect 320 -21 330 -17
rect 444 -24 448 -20
rect 546 -24 550 -20
rect 125 -38 129 -34
rect 302 -29 312 -25
rect 322 -29 332 -25
rect 347 -32 351 -28
rect 125 -46 129 -42
rect 161 -40 165 -36
rect 175 -40 179 -36
rect 193 -40 197 -36
rect 201 -40 205 -36
rect 109 -54 113 -50
rect 109 -62 113 -58
rect 109 -78 113 -74
rect 101 -85 105 -81
rect 355 -32 359 -28
rect 427 -32 431 -28
rect 435 -32 439 -28
rect 302 -37 314 -33
rect 320 -37 330 -33
rect 444 -40 448 -36
rect 546 -40 550 -36
rect 302 -45 312 -41
rect 322 -45 332 -41
rect 363 -48 367 -44
rect 395 -48 399 -44
rect 465 -48 469 -44
rect 161 -56 165 -52
rect 175 -56 179 -52
rect 193 -56 197 -52
rect 201 -56 205 -52
rect 302 -53 314 -49
rect 320 -53 330 -49
rect 444 -56 448 -52
rect 546 -56 550 -52
rect 125 -70 129 -66
rect 302 -61 312 -57
rect 322 -61 332 -57
rect 379 -64 383 -60
rect 395 -64 399 -60
rect 411 -64 415 -60
rect 481 -64 485 -60
rect 489 -64 493 -60
rect 125 -78 129 -74
rect 175 -72 179 -68
rect 193 -72 197 -68
rect 302 -69 314 -65
rect 320 -69 330 -65
rect 444 -72 448 -68
rect 546 -72 550 -68
rect 322 -77 332 -73
rect 117 -85 121 -81
rect 37 -110 41 -106
rect 45 -117 49 -113
rect 45 -133 49 -129
rect 45 -157 49 -153
rect 53 -110 57 -106
rect 69 -110 73 -106
rect 61 -157 65 -153
rect 45 -165 49 -161
rect 37 -172 41 -168
rect 53 -172 57 -168
rect 85 -110 89 -106
rect 77 -117 81 -113
rect 77 -125 81 -121
rect 77 -133 81 -129
rect 77 -141 81 -137
rect 77 -149 81 -145
rect 77 -165 81 -161
rect 69 -172 73 -168
rect 101 -110 105 -106
rect 117 -110 121 -106
rect 109 -117 113 -113
rect 109 -125 113 -121
rect 93 -133 97 -129
rect 93 -141 97 -137
rect 93 -149 97 -145
rect 93 -157 97 -153
rect 93 -165 97 -161
rect 85 -172 89 -168
rect 161 -103 165 -99
rect 201 -103 205 -99
rect 302 -108 312 -104
rect 363 -111 367 -107
rect 505 -80 509 -76
rect 161 -119 165 -115
rect 175 -119 179 -115
rect 193 -119 197 -115
rect 201 -119 205 -115
rect 302 -116 314 -112
rect 320 -116 330 -112
rect 444 -119 448 -115
rect 546 -119 550 -115
rect 125 -133 129 -129
rect 302 -124 312 -120
rect 322 -124 332 -120
rect 363 -127 367 -123
rect 387 -127 391 -123
rect 513 -127 517 -123
rect 125 -141 129 -137
rect 161 -135 165 -131
rect 175 -135 179 -131
rect 193 -135 197 -131
rect 201 -135 205 -131
rect 109 -149 113 -145
rect 109 -157 113 -153
rect 109 -165 113 -161
rect 101 -172 105 -168
rect 302 -132 314 -128
rect 320 -132 330 -128
rect 444 -135 448 -131
rect 546 -135 550 -131
rect 302 -140 312 -136
rect 322 -140 332 -136
rect 419 -143 423 -139
rect 521 -143 525 -139
rect 529 -143 533 -139
rect 125 -157 129 -153
rect 175 -151 179 -147
rect 193 -151 197 -147
rect 201 -151 205 -147
rect 302 -148 314 -144
rect 320 -148 330 -144
rect 444 -151 448 -147
rect 546 -151 550 -147
rect 125 -165 129 -161
rect 302 -156 312 -152
rect 322 -156 332 -152
rect 347 -159 351 -155
rect 117 -172 121 -168
rect 193 -167 197 -163
rect 363 -159 367 -155
rect 302 -164 314 -160
rect 444 -167 448 -163
rect 546 -167 550 -163
rect 35 -200 39 -187
rect 43 -198 47 -185
rect 27 -221 31 -208
rect 35 -221 39 -206
rect 51 -200 55 -187
rect 59 -198 63 -185
rect 43 -221 47 -208
rect 51 -221 55 -206
rect 67 -200 71 -187
rect 75 -198 79 -185
rect 59 -221 63 -208
rect 67 -221 71 -206
rect 83 -200 87 -187
rect 91 -198 95 -185
rect 75 -221 79 -208
rect 83 -221 87 -206
rect 99 -200 103 -187
rect 107 -198 111 -185
rect 91 -221 95 -208
rect 99 -221 103 -206
rect 115 -200 119 -187
rect 123 -198 127 -185
rect 363 -190 367 -181
rect 107 -221 111 -208
rect 115 -221 119 -206
rect 347 -208 351 -200
rect 123 -221 127 -208
rect 379 -190 383 -181
rect 363 -208 367 -200
rect 395 -190 399 -181
rect 379 -208 383 -200
rect 347 -360 351 -350
rect 41 -370 47 -366
rect 57 -370 63 -366
rect 73 -370 79 -366
rect 89 -370 95 -366
rect 105 -370 111 -366
rect 121 -370 127 -366
rect 411 -190 415 -181
rect 395 -208 399 -200
rect 363 -360 367 -350
rect 42 -383 46 -379
rect 58 -383 62 -379
rect 74 -383 78 -379
rect 90 -383 94 -379
rect 106 -383 110 -379
rect 427 -190 431 -181
rect 411 -208 415 -200
rect 379 -360 383 -350
rect 363 -379 367 -370
rect 443 -190 447 -181
rect 427 -208 431 -200
rect 395 -360 399 -350
rect 379 -379 383 -370
rect 481 -190 485 -181
rect 465 -208 469 -200
rect 411 -360 415 -350
rect 395 -379 399 -370
rect 497 -190 501 -181
rect 481 -208 485 -200
rect 427 -360 431 -350
rect 411 -379 415 -370
rect 513 -190 517 -181
rect 497 -208 501 -200
rect 465 -360 469 -350
rect 427 -379 431 -370
rect 529 -190 533 -181
rect 513 -208 517 -200
rect 481 -360 485 -350
rect 443 -379 447 -370
rect 545 -190 549 -181
rect 529 -208 533 -200
rect 497 -360 501 -350
rect 481 -379 485 -370
rect 513 -360 517 -350
rect 497 -379 501 -370
rect 529 -360 533 -350
rect 513 -379 517 -370
rect 529 -379 533 -370
rect 545 -379 549 -370
rect 122 -383 126 -379
<< pdcontact >>
rect 345 24 543 28
rect 347 16 351 20
rect 355 16 359 20
rect 363 16 367 20
rect 371 16 375 20
rect 379 16 383 20
rect 387 16 391 20
rect 395 16 399 20
rect 403 16 407 20
rect 411 16 415 20
rect 419 16 423 20
rect 427 16 431 20
rect 435 16 439 20
rect 465 16 469 20
rect 473 16 477 20
rect 481 16 485 20
rect 489 16 493 20
rect 497 16 501 20
rect 505 16 509 20
rect 513 16 517 20
rect 521 16 525 20
rect 529 16 533 20
rect 537 16 541 20
rect 143 8 149 12
rect 5 -80 9 0
rect 13 -6 17 -2
rect 13 -14 17 -10
rect 13 -22 17 -18
rect 13 -30 17 -26
rect 13 -38 17 -34
rect 13 -46 17 -42
rect 13 -54 17 -50
rect 13 -62 17 -58
rect 13 -70 17 -66
rect 13 -78 17 -74
rect 145 0 149 4
rect 217 8 223 12
rect 217 0 221 4
rect 275 3 290 7
rect 143 -8 149 -4
rect 145 -16 149 -12
rect 217 -8 223 -4
rect 242 -5 262 -1
rect 268 -5 290 -1
rect 217 -16 221 -12
rect 242 -13 260 -9
rect 275 -13 290 -9
rect 143 -24 149 -20
rect 145 -32 149 -28
rect 217 -24 223 -20
rect 242 -21 262 -17
rect 268 -21 290 -17
rect 217 -32 221 -28
rect 242 -29 260 -25
rect 275 -29 290 -25
rect 143 -40 149 -36
rect 145 -48 149 -44
rect 217 -40 223 -36
rect 242 -37 262 -33
rect 268 -37 290 -33
rect 217 -48 221 -44
rect 242 -45 260 -41
rect 275 -45 290 -41
rect 143 -56 149 -52
rect 145 -64 149 -60
rect 217 -56 223 -52
rect 242 -53 262 -49
rect 268 -53 290 -49
rect 217 -64 221 -60
rect 242 -61 260 -57
rect 275 -61 290 -57
rect 143 -72 149 -68
rect 217 -72 223 -68
rect 242 -69 262 -65
rect 268 -69 290 -65
rect 242 -77 260 -73
rect 5 -167 9 -111
rect 13 -117 17 -113
rect 13 -125 17 -121
rect 13 -133 17 -129
rect 13 -141 17 -137
rect 13 -149 17 -145
rect 13 -157 17 -153
rect 13 -165 17 -161
rect 143 -103 149 -99
rect 145 -111 149 -107
rect 217 -103 223 -99
rect 217 -111 221 -107
rect 275 -108 290 -104
rect 143 -119 149 -115
rect 145 -127 149 -123
rect 217 -119 223 -115
rect 242 -116 262 -112
rect 268 -116 290 -112
rect 217 -127 221 -123
rect 242 -124 260 -120
rect 275 -124 290 -120
rect 143 -135 149 -131
rect 145 -143 149 -139
rect 217 -135 223 -131
rect 242 -132 262 -128
rect 268 -132 290 -128
rect 217 -143 221 -139
rect 242 -140 260 -136
rect 275 -140 290 -136
rect 143 -151 149 -147
rect 217 -151 223 -147
rect 242 -148 262 -144
rect 268 -148 290 -144
rect 217 -159 221 -155
rect 242 -156 260 -152
rect 275 -156 290 -152
rect 217 -167 223 -163
rect 268 -164 290 -160
rect 27 -251 31 -233
rect 35 -260 39 -233
rect 35 -292 39 -266
rect 43 -251 47 -233
rect 43 -285 47 -266
rect 51 -260 55 -233
rect 51 -292 55 -266
rect 59 -251 63 -233
rect 59 -285 63 -266
rect 67 -260 71 -233
rect 67 -292 71 -266
rect 75 -251 79 -233
rect 75 -285 79 -266
rect 83 -260 87 -233
rect 83 -292 87 -266
rect 91 -251 95 -233
rect 91 -285 95 -266
rect 99 -260 103 -233
rect 99 -292 103 -266
rect 107 -251 111 -233
rect 107 -285 111 -266
rect 115 -260 119 -233
rect 115 -292 119 -266
rect 123 -251 127 -233
rect 347 -242 351 -220
rect 363 -242 367 -220
rect 123 -285 127 -266
rect 42 -309 46 -305
rect 58 -309 62 -305
rect 74 -309 78 -305
rect 90 -309 94 -305
rect 106 -309 110 -305
rect 122 -309 126 -305
rect 379 -242 383 -220
rect 363 -273 367 -252
rect 363 -312 367 -288
rect 41 -322 47 -318
rect 57 -322 63 -318
rect 73 -322 79 -318
rect 89 -322 95 -318
rect 105 -322 111 -318
rect 121 -322 127 -318
rect 42 -341 46 -337
rect 58 -341 62 -337
rect 74 -341 78 -337
rect 90 -341 94 -337
rect 106 -341 110 -337
rect 122 -341 126 -337
rect 347 -338 351 -316
rect 41 -354 47 -350
rect 57 -354 63 -350
rect 73 -354 79 -350
rect 89 -354 95 -350
rect 105 -354 111 -350
rect 121 -354 127 -350
rect 395 -242 399 -220
rect 379 -273 383 -252
rect 379 -312 383 -288
rect 363 -338 367 -316
rect 411 -242 415 -220
rect 395 -273 399 -252
rect 395 -312 399 -288
rect 379 -338 383 -316
rect 427 -242 431 -220
rect 411 -273 415 -252
rect 411 -312 415 -288
rect 395 -338 399 -316
rect 465 -242 469 -220
rect 427 -273 431 -252
rect 427 -312 431 -288
rect 411 -338 415 -316
rect 481 -242 485 -220
rect 443 -273 447 -252
rect 443 -312 447 -288
rect 427 -338 431 -316
rect 497 -242 501 -220
rect 481 -273 485 -252
rect 481 -312 485 -288
rect 465 -338 469 -316
rect 513 -242 517 -220
rect 497 -273 501 -252
rect 497 -312 501 -288
rect 481 -338 485 -316
rect 529 -242 533 -220
rect 513 -273 517 -252
rect 513 -312 517 -288
rect 497 -338 501 -316
rect 529 -273 533 -252
rect 529 -312 533 -288
rect 513 -338 517 -316
rect 545 -273 549 -252
rect 545 -312 549 -288
rect 529 -338 533 -316
<< psubstratepcontact >>
rect 29 26 129 30
rect 444 0 448 4
rect 546 0 550 4
rect 315 -5 319 -1
rect 444 -16 448 -12
rect 546 -16 550 -12
rect 315 -21 319 -17
rect 444 -32 448 -28
rect 546 -32 550 -28
rect 315 -37 319 -33
rect 444 -48 448 -44
rect 546 -48 550 -44
rect 315 -53 319 -49
rect 444 -64 448 -60
rect 546 -64 550 -60
rect 315 -69 319 -65
rect 29 -103 33 -99
rect 45 -103 49 -99
rect 61 -103 65 -99
rect 77 -103 81 -99
rect 93 -103 97 -99
rect 109 -103 113 -99
rect 320 -98 343 -94
rect 125 -103 129 -99
rect 444 -111 448 -76
rect 546 -111 550 -76
rect 315 -116 319 -112
rect 444 -127 448 -123
rect 546 -127 550 -123
rect 315 -132 319 -128
rect 444 -143 448 -139
rect 546 -143 550 -139
rect 315 -148 319 -144
rect 444 -159 448 -155
rect 546 -159 550 -155
rect 315 -164 319 -160
rect 315 -175 323 -171
rect 347 -180 351 -176
rect 363 -180 367 -176
rect 35 -205 39 -201
rect 51 -205 55 -201
rect 67 -205 71 -201
rect 83 -205 87 -201
rect 99 -205 103 -201
rect 379 -180 383 -176
rect 115 -205 119 -201
rect 395 -180 399 -176
rect 411 -180 415 -176
rect 32 -370 36 -366
rect 48 -370 52 -366
rect 64 -370 68 -366
rect 80 -370 84 -366
rect 96 -370 100 -366
rect 112 -370 116 -366
rect 128 -370 132 -366
rect 427 -180 431 -176
rect 443 -180 447 -176
rect 465 -180 469 -176
rect 481 -180 485 -176
rect 497 -180 501 -176
rect 513 -180 517 -176
rect 529 -180 533 -176
rect 545 -180 549 -176
rect 347 -384 351 -380
rect 363 -384 367 -380
rect 379 -384 383 -380
rect 395 -384 399 -380
rect 411 -384 415 -380
rect 427 -384 431 -380
rect 443 -384 447 -380
rect 465 -384 469 -380
rect 481 -384 485 -380
rect 497 -384 501 -380
rect 513 -384 517 -380
rect 529 -384 533 -380
rect 545 -384 549 -380
<< nsubstratencontact >>
rect 345 29 543 33
rect 138 8 142 12
rect 0 -80 4 0
rect 224 8 228 12
rect 138 -8 142 -4
rect 224 -8 228 -4
rect 263 -5 267 -1
rect 138 -24 142 -20
rect 224 -24 228 -20
rect 263 -21 267 -17
rect 138 -40 142 -36
rect 224 -40 228 -36
rect 263 -37 267 -33
rect 138 -56 142 -52
rect 224 -56 228 -52
rect 263 -53 267 -49
rect 138 -72 142 -68
rect 224 -72 228 -68
rect 263 -69 267 -65
rect 0 -167 4 -111
rect 138 -103 142 -99
rect 224 -103 228 -99
rect 138 -119 142 -115
rect 224 -119 228 -115
rect 263 -116 267 -112
rect 138 -135 142 -131
rect 224 -135 228 -131
rect 263 -132 267 -128
rect 138 -151 142 -147
rect 224 -151 228 -147
rect 263 -148 267 -144
rect 224 -167 228 -163
rect 263 -164 267 -160
rect 35 -265 39 -261
rect 51 -265 55 -261
rect 67 -265 71 -261
rect 83 -265 87 -261
rect 99 -265 103 -261
rect 115 -265 119 -261
rect 347 -278 351 -274
rect 363 -278 367 -274
rect 32 -322 36 -318
rect 48 -322 52 -318
rect 64 -322 68 -318
rect 80 -322 84 -318
rect 96 -322 100 -318
rect 112 -322 116 -318
rect 128 -322 132 -318
rect 32 -354 36 -350
rect 48 -354 52 -350
rect 64 -354 68 -350
rect 80 -354 84 -350
rect 96 -354 100 -350
rect 112 -354 116 -350
rect 128 -354 132 -350
rect 379 -278 383 -274
rect 395 -278 399 -274
rect 411 -278 415 -274
rect 444 -242 448 -220
rect 427 -278 431 -274
rect 443 -278 447 -274
rect 465 -278 469 -274
rect 481 -278 485 -274
rect 444 -338 448 -317
rect 497 -278 501 -274
rect 513 -278 517 -274
rect 529 -278 533 -274
rect 545 -278 549 -274
<< polysilicon >>
rect 340 21 347 23
rect 351 21 355 23
rect 359 21 363 23
rect 367 21 371 23
rect 375 21 379 23
rect 383 21 387 23
rect 391 21 395 23
rect 399 21 403 23
rect 407 21 411 23
rect 415 21 419 23
rect 423 21 427 23
rect 431 21 435 23
rect 439 21 465 23
rect 469 21 473 23
rect 477 21 481 23
rect 485 21 489 23
rect 493 21 497 23
rect 501 21 505 23
rect 509 21 513 23
rect 517 21 521 23
rect 525 21 529 23
rect 533 21 537 23
rect 541 21 548 23
rect 446 20 450 21
rect 10 -2 12 3
rect 10 -10 12 -6
rect 10 -18 12 -14
rect 10 -26 12 -22
rect 10 -34 12 -30
rect 10 -42 12 -38
rect 10 -50 12 -46
rect 10 -58 12 -54
rect 10 -66 12 -62
rect 10 -74 12 -70
rect 10 -87 12 -78
rect 34 -87 36 8
rect 42 -18 44 8
rect 42 -34 44 -22
rect 42 -50 44 -38
rect 42 -87 44 -54
rect 50 -87 52 8
rect 58 -87 60 8
rect 66 -87 68 8
rect 74 -87 76 8
rect 82 -66 84 8
rect 90 -2 92 8
rect 90 -26 92 -6
rect 90 -42 92 -30
rect 98 -34 100 8
rect 106 -2 108 8
rect 106 -10 108 -6
rect 114 -10 116 8
rect 122 -2 124 8
rect 143 5 145 7
rect 149 5 161 7
rect 165 5 168 7
rect 172 5 201 7
rect 205 5 217 7
rect 221 5 223 7
rect 135 -3 145 -1
rect 149 -3 172 -1
rect 176 -3 178 -1
rect 239 0 270 2
rect 290 0 302 2
rect 312 0 314 2
rect 190 -3 193 -1
rect 197 -3 217 -1
rect 221 -3 223 -1
rect 106 -18 108 -14
rect 114 -18 116 -14
rect 106 -26 108 -22
rect 114 -26 116 -22
rect 98 -42 100 -38
rect 90 -50 92 -46
rect 98 -50 100 -46
rect 90 -58 92 -54
rect 98 -58 100 -54
rect 82 -74 84 -70
rect 82 -87 84 -78
rect 90 -87 92 -62
rect 98 -87 100 -62
rect 106 -74 108 -30
rect 114 -50 116 -30
rect 122 -34 124 -6
rect 135 -12 137 -3
rect 143 -11 145 -9
rect 149 -11 161 -9
rect 165 -11 168 -9
rect 342 -3 371 -1
rect 375 -3 379 -1
rect 383 -3 451 -1
rect 239 -8 240 -6
rect 260 -8 322 -6
rect 332 -8 334 -6
rect 455 -3 537 -1
rect 541 -3 553 -1
rect 455 -5 460 -3
rect 172 -11 201 -9
rect 205 -11 217 -9
rect 221 -11 223 -9
rect 135 -19 145 -17
rect 149 -19 172 -17
rect 176 -19 178 -17
rect 342 -11 379 -9
rect 383 -11 451 -9
rect 239 -16 270 -14
rect 290 -16 302 -14
rect 312 -16 314 -14
rect 455 -11 553 -9
rect 190 -19 193 -17
rect 197 -19 217 -17
rect 221 -19 223 -17
rect 135 -28 137 -19
rect 143 -27 145 -25
rect 149 -27 161 -25
rect 165 -27 168 -25
rect 342 -19 355 -17
rect 359 -19 451 -17
rect 239 -24 240 -22
rect 260 -24 322 -22
rect 332 -24 334 -22
rect 455 -19 553 -17
rect 455 -21 460 -19
rect 172 -27 201 -25
rect 205 -27 217 -25
rect 221 -27 223 -25
rect 135 -35 145 -33
rect 149 -35 172 -33
rect 176 -35 178 -33
rect 342 -27 427 -25
rect 431 -27 435 -25
rect 439 -27 451 -25
rect 239 -32 270 -30
rect 290 -32 302 -30
rect 312 -32 314 -30
rect 190 -35 193 -33
rect 197 -35 217 -33
rect 221 -35 223 -33
rect 122 -42 124 -38
rect 135 -44 137 -35
rect 143 -43 145 -41
rect 149 -43 161 -41
rect 165 -43 168 -41
rect 114 -58 116 -54
rect 106 -87 108 -78
rect 114 -87 116 -62
rect 122 -66 124 -46
rect 455 -27 553 -25
rect 342 -35 347 -33
rect 351 -35 355 -33
rect 359 -35 451 -33
rect 239 -40 240 -38
rect 260 -40 322 -38
rect 332 -40 334 -38
rect 455 -35 553 -33
rect 455 -37 460 -35
rect 172 -43 201 -41
rect 205 -43 217 -41
rect 221 -43 223 -41
rect 135 -51 145 -49
rect 149 -51 172 -49
rect 176 -51 178 -49
rect 342 -43 395 -41
rect 399 -43 451 -41
rect 239 -48 270 -46
rect 290 -48 302 -46
rect 312 -48 314 -46
rect 455 -43 465 -41
rect 469 -43 553 -41
rect 455 -45 460 -43
rect 190 -51 193 -49
rect 197 -51 217 -49
rect 221 -51 223 -49
rect 135 -60 137 -51
rect 143 -59 145 -57
rect 149 -59 161 -57
rect 165 -59 168 -57
rect 342 -51 363 -49
rect 367 -51 451 -49
rect 239 -56 240 -54
rect 260 -56 322 -54
rect 332 -56 334 -54
rect 455 -51 553 -49
rect 455 -53 460 -51
rect 172 -59 201 -57
rect 205 -59 217 -57
rect 221 -59 223 -57
rect 135 -67 145 -65
rect 149 -67 172 -65
rect 176 -67 178 -65
rect 342 -59 379 -57
rect 383 -59 411 -57
rect 415 -59 451 -57
rect 239 -64 270 -62
rect 290 -64 302 -62
rect 312 -64 314 -62
rect 455 -59 481 -57
rect 485 -59 489 -57
rect 493 -59 553 -57
rect 455 -61 460 -59
rect 190 -67 193 -65
rect 197 -67 217 -65
rect 221 -67 223 -65
rect 122 -74 124 -70
rect 135 -76 137 -67
rect 342 -67 395 -65
rect 399 -67 451 -65
rect 239 -72 240 -70
rect 260 -72 322 -70
rect 332 -72 334 -70
rect 455 -67 553 -65
rect 455 -69 460 -67
rect 342 -75 451 -73
rect 122 -87 124 -78
rect 10 -113 12 -96
rect 10 -121 12 -117
rect 10 -129 12 -125
rect 10 -137 12 -133
rect 10 -145 12 -141
rect 10 -153 12 -149
rect 10 -161 12 -157
rect 10 -170 12 -165
rect 34 -175 36 -96
rect 42 -113 44 -96
rect 42 -129 44 -117
rect 42 -153 44 -133
rect 42 -161 44 -157
rect 50 -161 52 -96
rect 58 -153 60 -96
rect 66 -153 68 -96
rect 42 -175 44 -165
rect 50 -175 52 -165
rect 58 -175 60 -157
rect 66 -175 68 -157
rect 74 -161 76 -96
rect 82 -113 84 -96
rect 82 -121 84 -117
rect 82 -129 84 -125
rect 82 -137 84 -133
rect 82 -145 84 -141
rect 74 -175 76 -165
rect 82 -175 84 -149
rect 90 -153 92 -96
rect 98 -129 100 -96
rect 106 -113 108 -96
rect 114 -113 116 -96
rect 106 -121 108 -117
rect 114 -121 116 -117
rect 98 -137 100 -133
rect 98 -145 100 -141
rect 90 -161 92 -157
rect 90 -175 92 -165
rect 98 -175 100 -149
rect 106 -153 108 -125
rect 114 -145 116 -125
rect 122 -129 124 -96
rect 143 -106 145 -104
rect 149 -106 161 -104
rect 165 -106 168 -104
rect 172 -106 201 -104
rect 205 -106 217 -104
rect 221 -106 223 -104
rect 135 -114 145 -112
rect 149 -114 172 -112
rect 176 -114 178 -112
rect 239 -111 270 -109
rect 290 -111 302 -109
rect 312 -111 314 -109
rect 455 -75 505 -73
rect 509 -75 553 -73
rect 455 -77 460 -75
rect 190 -114 193 -112
rect 197 -114 217 -112
rect 221 -114 223 -112
rect 135 -123 137 -114
rect 143 -122 145 -120
rect 149 -122 161 -120
rect 165 -122 168 -120
rect 342 -114 363 -112
rect 367 -114 451 -112
rect 239 -119 240 -117
rect 260 -119 322 -117
rect 332 -119 334 -117
rect 455 -114 553 -112
rect 455 -116 460 -114
rect 172 -122 201 -120
rect 205 -122 217 -120
rect 221 -122 223 -120
rect 135 -130 145 -128
rect 149 -130 172 -128
rect 176 -130 178 -128
rect 342 -122 387 -120
rect 391 -122 451 -120
rect 239 -127 270 -125
rect 290 -127 302 -125
rect 312 -127 314 -125
rect 455 -122 513 -120
rect 517 -122 553 -120
rect 455 -124 460 -122
rect 190 -130 193 -128
rect 197 -130 217 -128
rect 221 -130 223 -128
rect 122 -137 124 -133
rect 135 -139 137 -130
rect 143 -138 145 -136
rect 149 -138 161 -136
rect 165 -138 168 -136
rect 106 -161 108 -157
rect 106 -175 108 -165
rect 114 -175 116 -149
rect 122 -153 124 -141
rect 342 -130 363 -128
rect 367 -130 451 -128
rect 239 -135 240 -133
rect 260 -135 322 -133
rect 332 -135 334 -133
rect 455 -130 553 -128
rect 455 -132 460 -130
rect 172 -138 201 -136
rect 205 -138 217 -136
rect 221 -138 223 -136
rect 135 -146 145 -144
rect 149 -146 172 -144
rect 176 -146 178 -144
rect 342 -138 451 -136
rect 239 -143 270 -141
rect 290 -143 302 -141
rect 312 -143 314 -141
rect 455 -138 521 -136
rect 525 -138 553 -136
rect 455 -140 460 -138
rect 190 -146 193 -144
rect 197 -146 217 -144
rect 221 -146 223 -144
rect 135 -155 137 -146
rect 342 -146 419 -144
rect 423 -146 451 -144
rect 239 -151 240 -149
rect 260 -151 322 -149
rect 332 -151 334 -149
rect 455 -146 529 -144
rect 533 -146 553 -144
rect 455 -148 460 -146
rect 172 -154 201 -152
rect 205 -154 217 -152
rect 221 -154 223 -152
rect 122 -161 124 -157
rect 342 -154 347 -152
rect 351 -154 451 -152
rect 239 -159 270 -157
rect 290 -159 302 -157
rect 312 -159 314 -157
rect 190 -162 193 -160
rect 197 -162 217 -160
rect 221 -162 223 -160
rect 122 -175 124 -165
rect 455 -154 553 -152
rect 342 -162 347 -160
rect 351 -162 363 -160
rect 367 -162 451 -160
rect 455 -162 553 -160
rect 455 -164 460 -162
rect 359 -173 362 -171
rect 375 -173 378 -171
rect 391 -173 394 -171
rect 407 -173 410 -171
rect 423 -173 426 -171
rect 439 -173 442 -171
rect 477 -173 480 -171
rect 493 -173 496 -171
rect 509 -173 512 -171
rect 525 -173 528 -171
rect 541 -173 544 -171
rect 360 -183 362 -173
rect 40 -185 42 -183
rect 56 -185 58 -183
rect 72 -185 74 -183
rect 88 -185 90 -183
rect 104 -185 106 -183
rect 120 -185 122 -183
rect 32 -208 34 -206
rect 32 -233 34 -221
rect 32 -295 34 -258
rect 40 -268 42 -198
rect 48 -208 50 -206
rect 48 -233 50 -221
rect 40 -295 42 -294
rect 48 -295 50 -258
rect 56 -268 58 -198
rect 64 -208 66 -206
rect 64 -233 66 -221
rect 56 -295 58 -294
rect 64 -295 66 -258
rect 72 -268 74 -198
rect 80 -208 82 -206
rect 80 -233 82 -221
rect 72 -295 74 -294
rect 80 -295 82 -258
rect 88 -268 90 -198
rect 96 -208 98 -206
rect 96 -233 98 -221
rect 88 -295 90 -294
rect 96 -295 98 -258
rect 104 -268 106 -198
rect 376 -183 378 -173
rect 352 -198 354 -197
rect 112 -208 114 -206
rect 112 -233 114 -221
rect 104 -295 106 -294
rect 112 -295 114 -258
rect 120 -268 122 -198
rect 352 -212 354 -208
rect 352 -220 354 -218
rect 352 -245 354 -244
rect 360 -247 362 -195
rect 392 -183 394 -173
rect 368 -198 370 -197
rect 368 -212 370 -208
rect 368 -220 370 -218
rect 368 -245 370 -244
rect 120 -295 122 -294
rect 39 -311 41 -310
rect 36 -312 41 -311
rect 45 -312 47 -310
rect 55 -311 57 -310
rect 52 -312 57 -311
rect 61 -312 63 -310
rect 71 -311 73 -310
rect 68 -312 73 -311
rect 77 -312 79 -310
rect 87 -311 89 -310
rect 84 -312 89 -311
rect 93 -312 95 -310
rect 103 -311 105 -310
rect 100 -312 105 -311
rect 109 -312 111 -310
rect 119 -311 121 -310
rect 116 -312 121 -311
rect 125 -312 127 -310
rect 38 -317 41 -315
rect 45 -317 47 -315
rect 54 -317 57 -315
rect 61 -317 63 -315
rect 70 -317 73 -315
rect 77 -317 79 -315
rect 86 -317 89 -315
rect 93 -317 95 -315
rect 102 -317 105 -315
rect 109 -317 111 -315
rect 118 -317 121 -315
rect 125 -317 127 -315
rect 352 -316 354 -249
rect 376 -247 378 -195
rect 408 -183 410 -173
rect 384 -198 386 -197
rect 384 -212 386 -208
rect 384 -220 386 -218
rect 384 -245 386 -244
rect 360 -273 362 -271
rect 360 -288 362 -285
rect 38 -325 40 -317
rect 54 -325 56 -317
rect 70 -325 72 -317
rect 86 -325 88 -317
rect 102 -325 104 -317
rect 118 -325 120 -317
rect 39 -343 41 -342
rect 36 -344 41 -343
rect 45 -344 47 -342
rect 55 -343 57 -342
rect 52 -344 57 -343
rect 61 -344 63 -342
rect 71 -343 73 -342
rect 68 -344 73 -343
rect 77 -344 79 -342
rect 87 -343 89 -342
rect 84 -344 89 -343
rect 93 -344 95 -342
rect 103 -343 105 -342
rect 100 -344 105 -343
rect 109 -344 111 -342
rect 352 -342 354 -338
rect 119 -343 121 -342
rect 116 -344 121 -343
rect 125 -344 127 -342
rect 38 -349 41 -347
rect 45 -349 47 -347
rect 54 -349 57 -347
rect 61 -349 63 -347
rect 70 -349 73 -347
rect 77 -349 79 -347
rect 86 -349 89 -347
rect 93 -349 95 -347
rect 102 -349 105 -347
rect 109 -349 111 -347
rect 118 -349 121 -347
rect 125 -349 127 -347
rect 38 -359 40 -349
rect 54 -359 56 -349
rect 70 -359 72 -349
rect 86 -359 88 -349
rect 102 -359 104 -349
rect 118 -359 120 -349
rect 352 -350 354 -348
rect 352 -363 354 -362
rect 38 -371 40 -363
rect 54 -371 56 -363
rect 70 -371 72 -363
rect 86 -371 88 -363
rect 102 -371 104 -363
rect 118 -371 120 -363
rect 360 -365 362 -312
rect 368 -316 370 -249
rect 392 -247 394 -195
rect 424 -183 426 -173
rect 400 -198 402 -197
rect 400 -212 402 -208
rect 400 -220 402 -218
rect 400 -245 402 -244
rect 376 -273 378 -271
rect 376 -288 378 -285
rect 368 -342 370 -338
rect 368 -350 370 -348
rect 368 -363 370 -362
rect 38 -373 41 -371
rect 45 -373 47 -371
rect 54 -373 57 -371
rect 61 -373 63 -371
rect 70 -373 73 -371
rect 77 -373 79 -371
rect 86 -373 89 -371
rect 93 -373 95 -371
rect 102 -373 105 -371
rect 109 -373 111 -371
rect 118 -373 121 -371
rect 125 -373 127 -371
rect 37 -377 41 -376
rect 39 -378 41 -377
rect 45 -378 47 -376
rect 53 -377 57 -376
rect 55 -378 57 -377
rect 61 -378 63 -376
rect 69 -377 73 -376
rect 71 -378 73 -377
rect 77 -378 79 -376
rect 85 -377 89 -376
rect 87 -378 89 -377
rect 93 -378 95 -376
rect 101 -377 105 -376
rect 103 -378 105 -377
rect 109 -378 111 -376
rect 117 -377 121 -376
rect 119 -378 121 -377
rect 125 -378 127 -376
rect 376 -365 378 -312
rect 384 -316 386 -249
rect 408 -247 410 -195
rect 440 -183 442 -173
rect 416 -198 418 -197
rect 416 -212 418 -208
rect 416 -220 418 -218
rect 416 -245 418 -244
rect 392 -273 394 -271
rect 392 -288 394 -285
rect 384 -342 386 -338
rect 384 -350 386 -348
rect 384 -363 386 -362
rect 360 -379 362 -377
rect 392 -365 394 -312
rect 400 -316 402 -249
rect 424 -247 426 -195
rect 478 -183 480 -173
rect 432 -198 434 -197
rect 432 -212 434 -208
rect 432 -220 434 -218
rect 432 -245 434 -244
rect 408 -273 410 -271
rect 408 -288 410 -285
rect 400 -342 402 -338
rect 400 -350 402 -348
rect 400 -363 402 -362
rect 376 -379 378 -377
rect 408 -365 410 -312
rect 416 -316 418 -249
rect 440 -247 442 -195
rect 494 -183 496 -173
rect 470 -198 472 -197
rect 470 -212 472 -208
rect 470 -220 472 -218
rect 470 -245 472 -244
rect 424 -273 426 -271
rect 424 -288 426 -285
rect 416 -342 418 -338
rect 416 -350 418 -348
rect 416 -363 418 -362
rect 392 -379 394 -377
rect 424 -365 426 -312
rect 432 -316 434 -249
rect 478 -247 480 -195
rect 510 -183 512 -173
rect 486 -198 488 -197
rect 486 -212 488 -208
rect 486 -220 488 -218
rect 486 -245 488 -244
rect 440 -273 442 -271
rect 440 -288 442 -285
rect 432 -342 434 -338
rect 432 -350 434 -348
rect 432 -363 434 -362
rect 408 -379 410 -377
rect 440 -365 442 -312
rect 470 -316 472 -249
rect 494 -247 496 -195
rect 526 -183 528 -173
rect 502 -198 504 -197
rect 502 -212 504 -208
rect 502 -220 504 -218
rect 502 -245 504 -244
rect 478 -273 480 -271
rect 478 -288 480 -285
rect 470 -342 472 -338
rect 470 -350 472 -348
rect 470 -363 472 -362
rect 424 -379 426 -377
rect 478 -365 480 -312
rect 486 -316 488 -249
rect 510 -247 512 -195
rect 542 -183 544 -173
rect 518 -198 520 -197
rect 518 -212 520 -208
rect 518 -220 520 -218
rect 518 -245 520 -244
rect 494 -273 496 -271
rect 494 -288 496 -285
rect 486 -342 488 -338
rect 486 -350 488 -348
rect 486 -363 488 -362
rect 440 -379 442 -377
rect 494 -365 496 -312
rect 502 -316 504 -249
rect 526 -247 528 -195
rect 534 -198 536 -197
rect 534 -212 536 -208
rect 534 -220 536 -218
rect 534 -245 536 -244
rect 510 -273 512 -271
rect 510 -288 512 -285
rect 502 -342 504 -338
rect 502 -350 504 -348
rect 502 -363 504 -362
rect 478 -379 480 -377
rect 510 -365 512 -312
rect 518 -316 520 -249
rect 542 -247 544 -195
rect 526 -273 528 -271
rect 526 -288 528 -285
rect 518 -342 520 -338
rect 518 -350 520 -348
rect 518 -363 520 -362
rect 494 -379 496 -377
rect 526 -365 528 -312
rect 534 -316 536 -249
rect 542 -273 544 -271
rect 542 -288 544 -285
rect 534 -342 536 -338
rect 534 -350 536 -348
rect 534 -363 536 -362
rect 510 -379 512 -377
rect 542 -365 544 -312
rect 526 -379 528 -377
rect 542 -379 544 -377
<< polycontact >>
rect 548 21 552 25
rect 338 17 342 21
rect 446 16 450 20
rect 34 8 38 12
rect 42 8 46 12
rect 50 8 54 12
rect 58 8 62 12
rect 66 8 70 12
rect 74 8 78 12
rect 82 8 86 12
rect 90 8 94 12
rect 98 8 102 12
rect 106 8 110 12
rect 114 8 118 12
rect 122 8 126 12
rect 8 3 12 7
rect 168 4 172 8
rect 186 -3 190 1
rect 235 -1 239 3
rect 131 -13 135 -9
rect 168 -12 172 -8
rect 338 -5 342 -1
rect 235 -9 239 -5
rect 451 -5 455 -1
rect 553 -5 557 -1
rect 186 -19 190 -15
rect 235 -17 239 -13
rect 338 -13 342 -9
rect 451 -13 455 -9
rect 553 -13 557 -9
rect 131 -29 135 -25
rect 168 -28 172 -24
rect 338 -21 342 -17
rect 235 -25 239 -21
rect 451 -21 455 -17
rect 553 -21 557 -17
rect 186 -35 190 -31
rect 235 -33 239 -29
rect 338 -29 342 -25
rect 131 -45 135 -41
rect 168 -44 172 -40
rect 451 -29 455 -25
rect 553 -29 557 -25
rect 338 -37 342 -33
rect 235 -41 239 -37
rect 451 -37 455 -33
rect 553 -37 557 -33
rect 186 -51 190 -47
rect 235 -49 239 -45
rect 338 -45 342 -41
rect 451 -45 455 -41
rect 553 -45 557 -41
rect 131 -61 135 -57
rect 168 -60 172 -56
rect 338 -53 342 -49
rect 235 -57 239 -53
rect 451 -53 455 -49
rect 553 -53 557 -49
rect 186 -67 190 -63
rect 235 -65 239 -61
rect 338 -61 342 -57
rect 451 -61 455 -57
rect 553 -61 557 -57
rect 131 -77 135 -73
rect 338 -69 342 -65
rect 235 -73 239 -69
rect 451 -69 455 -65
rect 553 -69 557 -65
rect 338 -77 342 -73
rect 8 -96 12 -92
rect 34 -96 38 -92
rect 42 -96 46 -92
rect 50 -96 54 -92
rect 58 -96 62 -92
rect 66 -96 70 -92
rect 74 -96 78 -92
rect 82 -96 86 -92
rect 90 -96 94 -92
rect 98 -96 102 -92
rect 106 -96 110 -92
rect 114 -96 118 -92
rect 122 -96 126 -92
rect 8 -174 12 -170
rect 168 -107 172 -103
rect 186 -114 190 -110
rect 235 -112 239 -108
rect 451 -77 455 -73
rect 553 -77 557 -73
rect 131 -124 135 -120
rect 168 -123 172 -119
rect 338 -116 342 -112
rect 235 -120 239 -116
rect 451 -116 455 -112
rect 553 -116 557 -112
rect 186 -130 190 -126
rect 235 -128 239 -124
rect 338 -124 342 -120
rect 451 -124 455 -120
rect 553 -124 557 -120
rect 131 -140 135 -136
rect 168 -139 172 -135
rect 338 -132 342 -128
rect 235 -136 239 -132
rect 451 -132 455 -128
rect 553 -132 557 -128
rect 186 -146 190 -142
rect 235 -144 239 -140
rect 338 -140 342 -136
rect 451 -140 455 -136
rect 553 -140 557 -136
rect 131 -156 135 -152
rect 168 -155 172 -151
rect 338 -148 342 -144
rect 235 -152 239 -148
rect 451 -148 455 -144
rect 553 -148 557 -144
rect 186 -162 190 -158
rect 235 -160 239 -156
rect 338 -156 342 -152
rect 451 -156 455 -152
rect 553 -156 557 -152
rect 338 -164 342 -160
rect 451 -164 455 -160
rect 553 -164 557 -160
rect 355 -173 359 -169
rect 371 -173 375 -169
rect 387 -173 391 -169
rect 403 -173 407 -169
rect 419 -173 423 -169
rect 435 -173 439 -169
rect 473 -173 477 -169
rect 489 -173 493 -169
rect 505 -173 509 -169
rect 521 -173 525 -169
rect 537 -173 541 -169
rect 34 -179 38 -175
rect 42 -179 46 -175
rect 50 -179 54 -175
rect 58 -179 62 -175
rect 66 -179 70 -175
rect 74 -179 78 -175
rect 82 -179 86 -175
rect 90 -179 94 -175
rect 98 -179 102 -175
rect 106 -179 110 -175
rect 114 -179 118 -175
rect 122 -179 126 -175
rect 351 -197 355 -193
rect 351 -249 355 -245
rect 367 -197 371 -193
rect 32 -299 36 -295
rect 40 -299 44 -295
rect 48 -299 52 -295
rect 56 -299 60 -295
rect 64 -299 68 -295
rect 72 -299 76 -295
rect 80 -299 84 -295
rect 88 -299 92 -295
rect 96 -299 100 -295
rect 104 -299 108 -295
rect 112 -299 116 -295
rect 120 -299 124 -295
rect 35 -311 39 -307
rect 51 -311 55 -307
rect 67 -311 71 -307
rect 83 -311 87 -307
rect 99 -311 103 -307
rect 115 -311 119 -307
rect 367 -249 371 -245
rect 383 -197 387 -193
rect 360 -285 364 -281
rect 37 -329 41 -325
rect 53 -329 57 -325
rect 69 -329 73 -325
rect 85 -329 89 -325
rect 101 -329 105 -325
rect 117 -329 121 -325
rect 35 -343 39 -339
rect 51 -343 55 -339
rect 67 -343 71 -339
rect 83 -343 87 -339
rect 99 -343 103 -339
rect 115 -343 119 -339
rect 37 -363 41 -359
rect 53 -363 57 -359
rect 69 -363 73 -359
rect 85 -363 89 -359
rect 101 -363 105 -359
rect 117 -363 121 -359
rect 351 -367 355 -363
rect 383 -249 387 -245
rect 399 -197 403 -193
rect 376 -285 380 -281
rect 35 -381 39 -377
rect 51 -381 55 -377
rect 67 -381 71 -377
rect 83 -381 87 -377
rect 99 -381 103 -377
rect 115 -381 119 -377
rect 367 -367 371 -363
rect 399 -249 403 -245
rect 415 -197 419 -193
rect 392 -285 396 -281
rect 383 -367 387 -363
rect 415 -249 419 -245
rect 431 -197 435 -193
rect 408 -285 412 -281
rect 399 -367 403 -363
rect 431 -249 435 -245
rect 469 -197 473 -193
rect 424 -285 428 -281
rect 415 -367 419 -363
rect 469 -249 473 -245
rect 485 -197 489 -193
rect 440 -285 444 -281
rect 431 -367 435 -363
rect 485 -249 489 -245
rect 501 -197 505 -193
rect 478 -285 482 -281
rect 469 -367 473 -363
rect 501 -249 505 -245
rect 517 -197 521 -193
rect 494 -285 498 -281
rect 485 -367 489 -363
rect 517 -249 521 -245
rect 533 -197 537 -193
rect 510 -285 514 -281
rect 501 -367 505 -363
rect 533 -249 537 -245
rect 526 -285 530 -281
rect 517 -367 521 -363
rect 542 -285 546 -281
rect 533 -367 537 -363
<< metal1 >>
rect 16 26 29 30
rect 129 26 319 32
rect 345 28 543 29
rect 16 24 129 26
rect 16 16 20 24
rect 142 8 143 12
rect 153 8 161 11
rect 169 8 172 12
rect 8 7 12 8
rect 30 2 37 5
rect 41 2 53 5
rect 57 2 69 5
rect 73 2 85 5
rect 89 2 101 5
rect 105 2 117 5
rect 121 2 125 5
rect 4 -80 5 0
rect 17 -6 93 -3
rect 97 -6 109 -3
rect 113 -6 125 -3
rect 129 -6 130 -2
rect 138 -4 142 8
rect 153 4 156 8
rect 149 1 152 4
rect 142 -8 143 -4
rect 153 -8 161 -5
rect 169 -8 172 4
rect 17 -14 109 -11
rect 129 -11 131 -10
rect 113 -13 131 -11
rect 113 -14 132 -13
rect 17 -22 45 -19
rect 49 -22 109 -19
rect 129 -19 130 -18
rect 113 -22 130 -19
rect 138 -20 142 -8
rect 153 -12 156 -8
rect 149 -15 152 -12
rect 142 -24 143 -20
rect 153 -24 161 -21
rect 169 -24 172 -12
rect 17 -30 93 -27
rect 97 -30 109 -27
rect 129 -27 131 -26
rect 113 -29 131 -27
rect 113 -30 132 -29
rect 17 -38 45 -35
rect 49 -38 93 -35
rect 97 -38 125 -35
rect 129 -38 130 -34
rect 138 -36 142 -24
rect 153 -28 156 -24
rect 149 -31 152 -28
rect 142 -40 143 -36
rect 153 -40 161 -37
rect 169 -40 172 -28
rect 17 -46 93 -43
rect 97 -46 125 -43
rect 129 -45 131 -42
rect 129 -46 132 -45
rect 17 -54 45 -51
rect 49 -54 93 -51
rect 97 -54 109 -51
rect 129 -51 130 -50
rect 113 -54 130 -51
rect 138 -52 142 -40
rect 153 -44 156 -40
rect 149 -47 152 -44
rect 142 -56 143 -52
rect 153 -56 161 -53
rect 169 -56 172 -44
rect 17 -62 93 -59
rect 97 -62 109 -59
rect 129 -59 131 -58
rect 113 -61 131 -59
rect 113 -62 132 -61
rect 17 -70 77 -67
rect 81 -70 125 -67
rect 129 -70 130 -66
rect 138 -68 142 -56
rect 153 -60 156 -56
rect 149 -63 152 -60
rect 142 -72 143 -68
rect 17 -78 77 -75
rect 81 -78 109 -75
rect 113 -78 125 -75
rect 129 -77 131 -74
rect 129 -78 132 -77
rect 1 -111 5 -80
rect 30 -84 37 -81
rect 41 -84 53 -81
rect 57 -84 69 -81
rect 73 -84 85 -81
rect 89 -84 101 -81
rect 105 -84 117 -81
rect 121 -84 125 -81
rect 138 -99 142 -72
rect 20 -103 29 -99
rect 33 -103 45 -99
rect 49 -103 61 -99
rect 65 -103 77 -99
rect 81 -103 93 -99
rect 97 -103 109 -99
rect 113 -103 125 -99
rect 142 -103 143 -99
rect 153 -103 161 -100
rect 169 -103 172 -60
rect 30 -109 37 -106
rect 41 -109 53 -106
rect 57 -109 69 -106
rect 73 -109 85 -106
rect 89 -109 101 -106
rect 105 -109 117 -106
rect 121 -109 125 -106
rect 4 -167 5 -111
rect 17 -117 45 -114
rect 49 -117 77 -114
rect 81 -117 109 -114
rect 129 -114 130 -113
rect 113 -117 130 -114
rect 138 -115 142 -103
rect 153 -107 156 -103
rect 149 -110 152 -107
rect 142 -119 143 -115
rect 153 -119 161 -116
rect 169 -119 172 -107
rect 17 -125 77 -122
rect 81 -125 109 -122
rect 129 -122 131 -121
rect 113 -124 131 -122
rect 113 -125 132 -124
rect 17 -133 45 -130
rect 49 -133 77 -130
rect 81 -133 93 -130
rect 97 -133 125 -130
rect 129 -133 130 -129
rect 138 -131 142 -119
rect 153 -123 156 -119
rect 149 -126 152 -123
rect 142 -135 143 -131
rect 153 -135 161 -132
rect 169 -135 172 -123
rect 17 -141 77 -138
rect 81 -141 93 -138
rect 97 -141 125 -138
rect 129 -140 131 -137
rect 129 -141 132 -140
rect 17 -149 77 -146
rect 81 -149 93 -146
rect 97 -149 109 -146
rect 129 -146 130 -145
rect 113 -149 130 -146
rect 138 -147 142 -135
rect 153 -139 156 -135
rect 149 -142 152 -139
rect 142 -151 143 -147
rect 169 -151 172 -139
rect 17 -157 45 -154
rect 49 -157 61 -154
rect 65 -157 93 -154
rect 97 -157 109 -154
rect 113 -157 125 -154
rect 129 -156 131 -153
rect 129 -157 132 -156
rect 17 -165 45 -162
rect 49 -165 77 -162
rect 81 -165 93 -162
rect 97 -165 109 -162
rect 113 -165 125 -162
rect 129 -165 130 -161
rect 138 -167 142 -151
rect 1 -288 5 -167
rect 30 -172 37 -169
rect 41 -172 53 -169
rect 57 -172 69 -169
rect 73 -172 85 -169
rect 89 -172 101 -169
rect 105 -172 117 -169
rect 121 -172 135 -169
rect 138 -171 147 -167
rect 8 -175 12 -174
rect 132 -179 135 -172
rect 1 -318 5 -292
rect 9 -310 12 -179
rect 35 -180 39 -179
rect 43 -180 47 -179
rect 51 -180 55 -179
rect 59 -180 63 -179
rect 67 -180 71 -179
rect 75 -180 79 -179
rect 83 -180 87 -179
rect 91 -180 95 -179
rect 99 -180 103 -179
rect 107 -180 111 -179
rect 115 -180 119 -179
rect 123 -180 127 -179
rect 43 -185 47 -184
rect 59 -185 63 -184
rect 35 -201 39 -200
rect 75 -185 79 -184
rect 51 -201 55 -200
rect 91 -185 95 -184
rect 67 -201 71 -200
rect 107 -185 111 -184
rect 83 -201 87 -200
rect 123 -185 127 -184
rect 99 -201 103 -200
rect 139 -187 147 -171
rect 169 -171 172 -155
rect 179 -179 183 26
rect 186 -4 190 -3
rect 193 -4 197 26
rect 224 15 308 19
rect 224 12 228 15
rect 205 8 211 11
rect 223 8 224 12
rect 208 4 211 8
rect 212 1 217 4
rect 224 -4 228 8
rect 268 -1 272 15
rect 315 10 319 26
rect 342 24 345 28
rect 543 24 545 28
rect 334 17 338 20
rect 548 20 552 21
rect 290 4 302 7
rect 293 -1 296 4
rect 315 6 338 10
rect 315 -1 319 6
rect 205 -8 211 -5
rect 223 -8 224 -4
rect 262 -5 263 -1
rect 267 -5 268 -1
rect 314 -5 315 -1
rect 319 -5 320 -1
rect 337 -5 338 -1
rect 186 -20 190 -19
rect 193 -20 197 -8
rect 208 -12 211 -8
rect 212 -15 217 -12
rect 224 -20 228 -8
rect 260 -13 261 -9
rect 268 -17 272 -5
rect 290 -12 302 -9
rect 293 -17 296 -12
rect 315 -17 319 -5
rect 332 -13 333 -9
rect 337 -13 338 -9
rect 205 -24 211 -21
rect 223 -24 224 -20
rect 262 -21 263 -17
rect 267 -21 268 -17
rect 314 -21 315 -17
rect 319 -21 320 -17
rect 337 -21 338 -17
rect 186 -36 190 -35
rect 193 -36 197 -24
rect 208 -28 211 -24
rect 212 -31 217 -28
rect 224 -36 228 -24
rect 260 -29 261 -25
rect 268 -33 272 -21
rect 290 -28 302 -25
rect 293 -33 296 -28
rect 315 -33 319 -21
rect 332 -29 333 -25
rect 337 -29 338 -25
rect 347 -28 350 16
rect 355 -12 358 16
rect 355 -28 358 -16
rect 205 -40 211 -37
rect 223 -40 224 -36
rect 262 -37 263 -33
rect 267 -37 268 -33
rect 314 -37 315 -33
rect 319 -37 320 -33
rect 337 -37 338 -33
rect 186 -52 190 -51
rect 193 -52 197 -40
rect 208 -44 211 -40
rect 212 -47 217 -44
rect 224 -52 228 -40
rect 260 -45 261 -41
rect 268 -49 272 -37
rect 290 -44 302 -41
rect 293 -49 296 -44
rect 315 -49 319 -37
rect 332 -45 333 -41
rect 337 -45 338 -41
rect 205 -56 211 -53
rect 223 -56 224 -52
rect 262 -53 263 -49
rect 267 -53 268 -49
rect 314 -53 315 -49
rect 319 -53 320 -49
rect 337 -53 338 -49
rect 186 -68 190 -67
rect 193 -68 197 -56
rect 208 -60 211 -56
rect 212 -63 217 -60
rect 224 -68 228 -56
rect 260 -61 261 -57
rect 268 -65 272 -53
rect 290 -60 302 -57
rect 293 -65 296 -60
rect 315 -65 319 -53
rect 332 -61 333 -57
rect 337 -61 338 -57
rect 223 -72 224 -68
rect 262 -69 263 -65
rect 267 -69 268 -65
rect 314 -69 315 -65
rect 319 -69 320 -65
rect 337 -69 338 -65
rect 186 -115 190 -114
rect 193 -115 197 -72
rect 224 -99 228 -72
rect 260 -77 261 -73
rect 205 -103 211 -100
rect 223 -103 224 -99
rect 208 -107 211 -103
rect 212 -110 217 -107
rect 224 -115 228 -103
rect 268 -112 272 -69
rect 315 -94 319 -69
rect 332 -77 333 -73
rect 337 -77 338 -73
rect 319 -98 320 -94
rect 290 -107 302 -104
rect 293 -112 296 -107
rect 315 -112 319 -98
rect 205 -119 211 -116
rect 223 -119 224 -115
rect 262 -116 263 -112
rect 267 -116 268 -112
rect 314 -116 315 -112
rect 319 -116 320 -112
rect 337 -116 338 -112
rect 186 -131 190 -130
rect 193 -131 197 -119
rect 208 -123 211 -119
rect 212 -126 217 -123
rect 224 -131 228 -119
rect 260 -124 261 -120
rect 268 -128 272 -116
rect 290 -123 302 -120
rect 293 -128 296 -123
rect 315 -128 319 -116
rect 332 -124 333 -120
rect 337 -124 338 -120
rect 205 -135 211 -132
rect 223 -135 224 -131
rect 262 -132 263 -128
rect 267 -132 268 -128
rect 314 -132 315 -128
rect 319 -132 320 -128
rect 337 -132 338 -128
rect 186 -147 190 -146
rect 193 -147 197 -135
rect 208 -139 211 -135
rect 212 -142 217 -139
rect 224 -147 228 -135
rect 260 -140 261 -136
rect 268 -144 272 -132
rect 290 -139 302 -136
rect 293 -144 296 -139
rect 315 -144 319 -132
rect 332 -140 333 -136
rect 337 -140 338 -136
rect 205 -151 211 -148
rect 223 -151 224 -147
rect 262 -148 263 -144
rect 267 -148 268 -144
rect 314 -148 315 -144
rect 319 -148 320 -144
rect 337 -148 338 -144
rect 186 -163 190 -162
rect 193 -163 197 -151
rect 208 -155 211 -151
rect 212 -158 217 -155
rect 224 -163 228 -151
rect 260 -156 261 -152
rect 268 -160 272 -148
rect 290 -155 302 -152
rect 293 -160 296 -155
rect 315 -160 319 -148
rect 332 -156 333 -152
rect 337 -156 338 -152
rect 347 -155 350 -32
rect 223 -167 224 -163
rect 267 -164 268 -160
rect 314 -164 315 -160
rect 337 -164 338 -160
rect 139 -191 143 -187
rect 115 -201 119 -200
rect 9 -342 12 -314
rect 20 -205 35 -201
rect 39 -205 51 -201
rect 55 -205 67 -201
rect 71 -205 83 -201
rect 87 -205 99 -201
rect 103 -205 115 -201
rect 119 -205 132 -201
rect 16 -366 20 -205
rect 35 -206 39 -205
rect 51 -206 55 -205
rect 67 -206 71 -205
rect 83 -206 87 -205
rect 99 -206 103 -205
rect 115 -206 119 -205
rect 27 -226 30 -221
rect 27 -229 35 -226
rect 43 -226 46 -221
rect 43 -229 51 -226
rect 59 -226 62 -221
rect 59 -229 67 -226
rect 75 -226 78 -221
rect 75 -229 83 -226
rect 91 -226 94 -221
rect 91 -229 99 -226
rect 107 -226 110 -221
rect 107 -229 115 -226
rect 27 -233 30 -229
rect 43 -233 46 -229
rect 59 -233 62 -229
rect 75 -233 78 -229
rect 91 -233 94 -229
rect 107 -233 110 -229
rect 123 -233 126 -221
rect 29 -258 35 -254
rect 39 -258 51 -254
rect 35 -261 39 -260
rect 55 -258 67 -254
rect 51 -261 55 -260
rect 71 -258 83 -254
rect 67 -261 71 -260
rect 87 -258 99 -254
rect 83 -261 87 -260
rect 103 -258 115 -254
rect 99 -261 103 -260
rect 139 -254 147 -191
rect 119 -258 147 -254
rect 115 -261 119 -260
rect 35 -266 39 -265
rect 29 -292 35 -288
rect 43 -266 47 -265
rect 51 -266 55 -265
rect 39 -292 51 -288
rect 59 -266 63 -265
rect 67 -266 71 -265
rect 55 -292 67 -288
rect 75 -266 79 -265
rect 83 -266 87 -265
rect 71 -292 83 -288
rect 91 -266 95 -265
rect 99 -266 103 -265
rect 87 -292 99 -288
rect 107 -266 111 -265
rect 115 -266 119 -265
rect 103 -292 115 -288
rect 123 -266 127 -265
rect 139 -288 147 -258
rect 119 -292 143 -288
rect 33 -300 37 -299
rect 41 -300 45 -299
rect 49 -300 53 -299
rect 57 -300 61 -299
rect 65 -300 69 -299
rect 73 -300 77 -299
rect 81 -300 85 -299
rect 89 -300 93 -299
rect 97 -300 101 -299
rect 105 -300 109 -299
rect 113 -300 117 -299
rect 121 -300 125 -299
rect 42 -305 45 -304
rect 58 -305 61 -304
rect 74 -305 77 -304
rect 90 -305 93 -304
rect 106 -305 109 -304
rect 122 -305 125 -304
rect 35 -312 39 -311
rect 51 -312 55 -311
rect 67 -312 71 -311
rect 83 -312 87 -311
rect 99 -312 103 -311
rect 115 -312 119 -311
rect 29 -314 132 -312
rect 26 -315 132 -314
rect 139 -318 147 -292
rect 29 -322 32 -318
rect 36 -322 41 -318
rect 47 -322 48 -318
rect 52 -322 57 -318
rect 63 -322 64 -318
rect 68 -322 73 -318
rect 79 -322 80 -318
rect 84 -322 89 -318
rect 95 -322 96 -318
rect 100 -322 105 -318
rect 111 -322 112 -318
rect 116 -322 121 -318
rect 127 -322 128 -318
rect 132 -322 147 -318
rect 41 -329 42 -325
rect 57 -329 58 -325
rect 73 -329 74 -325
rect 89 -329 90 -325
rect 105 -329 106 -325
rect 121 -329 122 -325
rect 38 -336 45 -333
rect 54 -336 61 -333
rect 70 -336 77 -333
rect 86 -336 93 -333
rect 102 -336 109 -333
rect 118 -336 125 -333
rect 42 -337 45 -336
rect 58 -337 61 -336
rect 74 -337 77 -336
rect 90 -337 93 -336
rect 106 -337 109 -336
rect 122 -337 125 -336
rect 35 -344 39 -343
rect 51 -344 55 -343
rect 67 -344 71 -343
rect 83 -344 87 -343
rect 99 -344 103 -343
rect 115 -344 119 -343
rect 29 -346 132 -344
rect 26 -347 132 -346
rect 139 -350 147 -322
rect 29 -354 32 -350
rect 36 -354 41 -350
rect 47 -354 48 -350
rect 52 -354 57 -350
rect 63 -354 64 -350
rect 68 -354 73 -350
rect 79 -354 80 -350
rect 84 -354 89 -350
rect 95 -354 96 -350
rect 100 -354 105 -350
rect 111 -354 112 -350
rect 116 -354 121 -350
rect 127 -354 128 -350
rect 132 -354 147 -350
rect 41 -363 42 -359
rect 57 -363 58 -359
rect 73 -363 74 -359
rect 89 -363 90 -359
rect 105 -363 106 -359
rect 121 -363 122 -359
rect 16 -370 32 -366
rect 36 -370 41 -366
rect 47 -370 48 -366
rect 52 -370 57 -366
rect 63 -370 64 -366
rect 68 -370 73 -366
rect 79 -370 80 -366
rect 84 -370 89 -366
rect 95 -370 96 -366
rect 100 -370 105 -366
rect 111 -370 112 -366
rect 116 -370 121 -366
rect 127 -370 128 -366
rect 29 -376 132 -373
rect 35 -377 39 -376
rect 51 -377 55 -376
rect 67 -377 71 -376
rect 83 -377 87 -376
rect 99 -377 103 -376
rect 115 -377 119 -376
rect 42 -384 45 -383
rect 58 -384 61 -383
rect 74 -384 77 -383
rect 90 -384 93 -383
rect 106 -384 109 -383
rect 122 -384 125 -383
rect 38 -387 45 -384
rect 54 -387 61 -384
rect 70 -387 77 -384
rect 86 -387 93 -384
rect 102 -387 109 -384
rect 118 -387 125 -384
rect 139 -387 147 -354
rect 193 -179 197 -167
rect 151 -373 154 -183
rect 179 -201 183 -183
rect 224 -187 228 -167
rect 268 -187 272 -164
rect 315 -167 319 -164
rect 347 -167 350 -159
rect 355 -167 358 -32
rect 363 -44 366 16
rect 371 4 374 16
rect 379 4 382 16
rect 363 -107 366 -48
rect 363 -123 366 -111
rect 363 -155 366 -127
rect 363 -167 366 -159
rect 371 -167 374 0
rect 379 -12 382 0
rect 379 -60 382 -16
rect 379 -167 382 -64
rect 387 -123 390 16
rect 395 -44 398 16
rect 395 -60 398 -48
rect 387 -167 390 -127
rect 395 -167 398 -64
rect 403 -167 406 16
rect 411 -60 414 16
rect 411 -167 414 -64
rect 419 -139 422 16
rect 427 -28 430 16
rect 435 -28 438 16
rect 444 4 448 6
rect 444 -4 448 0
rect 444 -12 448 -8
rect 444 -20 448 -16
rect 444 -28 448 -24
rect 419 -167 422 -143
rect 427 -167 430 -32
rect 435 -167 438 -32
rect 444 -36 448 -32
rect 444 -44 448 -40
rect 465 -44 468 16
rect 444 -52 448 -48
rect 444 -60 448 -56
rect 444 -68 448 -64
rect 444 -76 448 -72
rect 448 -98 449 -94
rect 444 -115 448 -111
rect 444 -123 448 -119
rect 444 -131 448 -127
rect 444 -139 448 -135
rect 444 -147 448 -143
rect 444 -155 448 -151
rect 444 -163 448 -159
rect 465 -167 468 -48
rect 473 -167 476 16
rect 481 -60 484 16
rect 489 -60 492 16
rect 481 -167 484 -64
rect 489 -167 492 -64
rect 497 -167 500 16
rect 505 -76 508 16
rect 505 -167 508 -80
rect 513 -123 516 16
rect 513 -167 516 -127
rect 521 -139 524 16
rect 529 -139 532 16
rect 537 4 540 16
rect 546 4 550 6
rect 521 -167 524 -143
rect 529 -167 532 -143
rect 537 -167 540 0
rect 546 -4 550 0
rect 557 -5 558 -1
rect 546 -12 550 -8
rect 557 -13 558 -9
rect 546 -20 550 -16
rect 557 -21 558 -17
rect 546 -28 550 -24
rect 557 -29 558 -25
rect 546 -36 550 -32
rect 557 -37 558 -33
rect 546 -44 550 -40
rect 557 -45 558 -41
rect 546 -52 550 -48
rect 557 -53 558 -49
rect 546 -60 550 -56
rect 557 -61 558 -57
rect 546 -68 550 -64
rect 557 -69 558 -65
rect 546 -76 550 -72
rect 557 -77 558 -73
rect 550 -98 551 -94
rect 546 -115 550 -111
rect 557 -116 558 -112
rect 546 -123 550 -119
rect 557 -124 558 -120
rect 546 -131 550 -127
rect 557 -132 558 -128
rect 546 -139 550 -135
rect 557 -140 558 -136
rect 546 -147 550 -143
rect 557 -148 558 -144
rect 546 -155 550 -151
rect 557 -156 558 -152
rect 546 -163 550 -159
rect 557 -164 558 -160
rect 315 -171 323 -167
rect 347 -169 351 -167
rect 355 -169 359 -167
rect 363 -169 367 -167
rect 371 -169 375 -167
rect 379 -169 383 -167
rect 387 -169 391 -167
rect 395 -169 399 -167
rect 403 -169 407 -167
rect 411 -169 415 -167
rect 419 -169 423 -167
rect 427 -169 431 -167
rect 435 -169 439 -167
rect 465 -169 469 -167
rect 473 -169 477 -167
rect 481 -169 485 -167
rect 489 -169 493 -167
rect 497 -169 501 -167
rect 505 -169 509 -167
rect 513 -169 517 -167
rect 521 -169 525 -167
rect 529 -169 533 -167
rect 537 -169 541 -167
rect 308 -193 311 -175
rect 315 -176 323 -175
rect 315 -179 347 -176
rect 319 -180 347 -179
rect 351 -180 363 -176
rect 367 -180 379 -176
rect 383 -180 395 -176
rect 399 -180 411 -176
rect 415 -180 427 -176
rect 431 -180 443 -176
rect 447 -180 465 -176
rect 469 -180 481 -176
rect 485 -180 497 -176
rect 501 -180 513 -176
rect 517 -180 529 -176
rect 533 -180 545 -176
rect 319 -183 323 -180
rect 159 -343 162 -315
rect 151 -387 154 -377
rect 159 -387 162 -347
rect 300 -384 303 -249
rect 308 -364 311 -197
rect 308 -384 311 -368
rect 315 -380 323 -183
rect 363 -181 367 -180
rect 379 -181 383 -180
rect 395 -181 399 -180
rect 411 -181 415 -180
rect 427 -181 431 -180
rect 443 -181 447 -180
rect 481 -181 485 -180
rect 497 -181 501 -180
rect 513 -181 517 -180
rect 529 -181 533 -180
rect 545 -181 549 -180
rect 343 -197 351 -194
rect 355 -197 367 -194
rect 371 -197 383 -194
rect 387 -197 399 -194
rect 403 -197 415 -194
rect 419 -197 431 -194
rect 435 -197 469 -194
rect 473 -197 485 -194
rect 489 -197 501 -194
rect 505 -197 517 -194
rect 521 -197 533 -194
rect 537 -197 549 -194
rect 347 -213 350 -208
rect 363 -213 366 -208
rect 379 -213 382 -208
rect 395 -213 398 -208
rect 411 -213 414 -208
rect 427 -213 430 -208
rect 465 -213 468 -208
rect 481 -213 484 -208
rect 497 -213 500 -208
rect 513 -213 516 -208
rect 529 -213 532 -208
rect 347 -220 350 -217
rect 363 -220 366 -217
rect 379 -220 382 -217
rect 395 -220 398 -217
rect 411 -220 414 -217
rect 427 -220 430 -217
rect 444 -220 448 -219
rect 465 -220 468 -217
rect 481 -220 484 -217
rect 497 -220 500 -217
rect 513 -220 516 -217
rect 529 -220 532 -217
rect 343 -249 351 -246
rect 355 -249 367 -246
rect 371 -249 383 -246
rect 387 -249 399 -246
rect 403 -249 415 -246
rect 419 -249 431 -246
rect 435 -249 469 -246
rect 473 -249 485 -246
rect 489 -249 501 -246
rect 505 -249 517 -246
rect 521 -249 533 -246
rect 537 -249 549 -246
rect 363 -274 367 -273
rect 379 -274 383 -273
rect 395 -274 399 -273
rect 411 -274 415 -273
rect 427 -274 431 -273
rect 443 -274 447 -273
rect 481 -274 485 -273
rect 497 -274 501 -273
rect 513 -274 517 -273
rect 529 -274 533 -273
rect 545 -274 549 -273
rect 339 -278 347 -274
rect 351 -278 363 -274
rect 367 -278 379 -274
rect 383 -278 395 -274
rect 399 -278 411 -274
rect 415 -278 427 -274
rect 431 -278 443 -274
rect 447 -278 465 -274
rect 469 -278 481 -274
rect 485 -278 497 -274
rect 501 -278 513 -274
rect 517 -278 529 -274
rect 533 -278 545 -274
rect 339 -288 343 -278
rect 359 -285 360 -281
rect 375 -285 376 -281
rect 391 -285 392 -281
rect 407 -285 408 -281
rect 423 -285 424 -281
rect 439 -285 440 -281
rect 477 -285 478 -281
rect 493 -285 494 -281
rect 509 -285 510 -281
rect 525 -285 526 -281
rect 541 -285 542 -281
rect 343 -292 363 -288
rect 367 -292 379 -288
rect 383 -292 395 -288
rect 399 -292 411 -288
rect 415 -292 427 -288
rect 431 -292 443 -288
rect 447 -292 481 -288
rect 447 -312 448 -292
rect 485 -292 497 -288
rect 501 -292 513 -288
rect 517 -292 529 -288
rect 533 -292 545 -288
rect 444 -317 448 -312
rect 347 -343 350 -338
rect 363 -343 366 -338
rect 379 -343 382 -338
rect 395 -343 398 -338
rect 411 -343 414 -338
rect 427 -343 430 -338
rect 444 -343 448 -338
rect 465 -343 468 -338
rect 481 -343 484 -338
rect 497 -343 500 -338
rect 513 -343 516 -338
rect 529 -343 532 -338
rect 347 -350 350 -347
rect 363 -350 366 -347
rect 379 -350 382 -347
rect 395 -350 398 -347
rect 411 -350 414 -347
rect 427 -350 430 -347
rect 465 -350 468 -347
rect 481 -350 484 -347
rect 497 -350 500 -347
rect 513 -350 516 -347
rect 529 -350 532 -347
rect 343 -367 351 -364
rect 355 -367 367 -364
rect 371 -367 383 -364
rect 387 -367 399 -364
rect 403 -367 415 -364
rect 419 -367 431 -364
rect 435 -367 469 -364
rect 473 -367 485 -364
rect 489 -367 501 -364
rect 505 -367 517 -364
rect 521 -367 533 -364
rect 537 -367 549 -364
rect 363 -380 367 -379
rect 379 -380 383 -379
rect 395 -380 399 -379
rect 411 -380 415 -379
rect 427 -380 431 -379
rect 443 -380 447 -379
rect 481 -380 485 -379
rect 497 -380 501 -379
rect 513 -380 517 -379
rect 529 -380 533 -379
rect 545 -380 549 -379
rect 315 -384 347 -380
rect 351 -384 363 -380
rect 367 -384 379 -380
rect 383 -384 395 -380
rect 399 -384 411 -380
rect 415 -384 427 -380
rect 431 -384 443 -380
rect 447 -384 465 -380
rect 469 -384 481 -380
rect 485 -384 497 -380
rect 501 -384 513 -380
rect 517 -384 529 -380
rect 533 -384 545 -380
<< m2contact >>
rect 16 12 20 16
rect 34 12 38 16
rect 8 8 12 12
rect 42 12 46 16
rect 50 12 54 16
rect 58 12 62 16
rect 66 12 70 16
rect 74 12 78 16
rect 82 12 86 16
rect 90 12 94 16
rect 98 12 102 16
rect 106 12 110 16
rect 114 12 118 16
rect 122 12 126 16
rect 26 1 30 5
rect 130 -6 134 -2
rect 152 0 156 4
rect 130 -22 134 -18
rect 152 -16 156 -12
rect 130 -38 134 -34
rect 152 -32 156 -28
rect 130 -54 134 -50
rect 152 -48 156 -44
rect 130 -70 134 -66
rect 152 -64 156 -60
rect 26 -85 30 -81
rect 8 -92 12 -88
rect 34 -92 38 -88
rect 42 -92 46 -88
rect 50 -92 54 -88
rect 58 -92 62 -88
rect 66 -92 70 -88
rect 74 -92 78 -88
rect 82 -92 86 -88
rect 90 -92 94 -88
rect 98 -92 102 -88
rect 106 -92 110 -88
rect 114 -92 118 -88
rect 122 -92 126 -88
rect 16 -103 20 -99
rect 26 -110 30 -106
rect 130 -117 134 -113
rect 152 -111 156 -107
rect 130 -133 134 -129
rect 152 -127 156 -123
rect 130 -149 134 -145
rect 152 -143 156 -139
rect 130 -165 134 -161
rect 26 -172 30 -168
rect 8 -179 12 -175
rect 1 -292 5 -288
rect 35 -184 39 -180
rect 43 -184 47 -180
rect 51 -184 55 -180
rect 59 -184 63 -180
rect 67 -184 71 -180
rect 75 -184 79 -180
rect 83 -184 87 -180
rect 91 -184 95 -180
rect 99 -184 103 -180
rect 107 -184 111 -180
rect 115 -184 119 -180
rect 123 -184 127 -180
rect 132 -183 136 -179
rect 169 -175 173 -171
rect 186 -8 190 -4
rect 308 15 312 19
rect 208 0 212 4
rect 231 -1 235 3
rect 338 24 342 28
rect 330 16 334 20
rect 442 16 446 20
rect 548 16 552 20
rect 338 6 342 10
rect 293 -5 297 -1
rect 333 -5 337 -1
rect 186 -24 190 -20
rect 208 -16 212 -12
rect 231 -9 235 -5
rect 261 -13 265 -9
rect 231 -17 235 -13
rect 333 -13 337 -9
rect 293 -21 297 -17
rect 333 -21 337 -17
rect 186 -40 190 -36
rect 208 -32 212 -28
rect 231 -25 235 -21
rect 261 -29 265 -25
rect 231 -33 235 -29
rect 333 -29 337 -25
rect 293 -37 297 -33
rect 333 -37 337 -33
rect 186 -56 190 -52
rect 208 -48 212 -44
rect 231 -41 235 -37
rect 261 -45 265 -41
rect 231 -49 235 -45
rect 333 -45 337 -41
rect 293 -53 297 -49
rect 333 -53 337 -49
rect 186 -72 190 -68
rect 208 -64 212 -60
rect 231 -57 235 -53
rect 261 -61 265 -57
rect 231 -65 235 -61
rect 333 -61 337 -57
rect 293 -69 297 -65
rect 333 -69 337 -65
rect 186 -119 190 -115
rect 231 -73 235 -69
rect 261 -77 265 -73
rect 208 -111 212 -107
rect 231 -112 235 -108
rect 333 -77 337 -73
rect 315 -98 319 -94
rect 293 -116 297 -112
rect 333 -116 337 -112
rect 186 -135 190 -131
rect 208 -127 212 -123
rect 231 -120 235 -116
rect 261 -124 265 -120
rect 231 -128 235 -124
rect 333 -124 337 -120
rect 293 -132 297 -128
rect 333 -132 337 -128
rect 186 -151 190 -147
rect 208 -143 212 -139
rect 231 -136 235 -132
rect 261 -140 265 -136
rect 231 -144 235 -140
rect 333 -140 337 -136
rect 293 -148 297 -144
rect 333 -148 337 -144
rect 186 -167 190 -163
rect 208 -159 212 -155
rect 231 -152 235 -148
rect 261 -156 265 -152
rect 231 -160 235 -156
rect 333 -156 337 -152
rect 293 -164 297 -160
rect 333 -164 337 -160
rect 143 -191 147 -187
rect 8 -314 12 -310
rect 1 -322 5 -318
rect 8 -346 12 -342
rect 16 -205 20 -201
rect 132 -205 136 -201
rect 35 -229 39 -225
rect 51 -229 55 -225
rect 67 -229 71 -225
rect 83 -229 87 -225
rect 99 -229 103 -225
rect 115 -229 119 -225
rect 25 -292 29 -288
rect 43 -265 47 -261
rect 59 -265 63 -261
rect 75 -265 79 -261
rect 91 -265 95 -261
rect 107 -265 111 -261
rect 123 -265 127 -261
rect 143 -292 147 -288
rect 33 -304 37 -300
rect 41 -304 45 -300
rect 49 -304 53 -300
rect 57 -304 61 -300
rect 65 -304 69 -300
rect 73 -304 77 -300
rect 81 -304 85 -300
rect 89 -304 93 -300
rect 97 -304 101 -300
rect 105 -304 109 -300
rect 113 -304 117 -300
rect 121 -304 125 -300
rect 25 -314 29 -310
rect 132 -315 136 -311
rect 25 -322 29 -318
rect 42 -329 46 -325
rect 58 -329 62 -325
rect 74 -329 78 -325
rect 90 -329 94 -325
rect 106 -329 110 -325
rect 122 -329 126 -325
rect 34 -336 38 -332
rect 50 -336 54 -332
rect 66 -336 70 -332
rect 82 -336 86 -332
rect 98 -336 102 -332
rect 114 -336 118 -332
rect 25 -346 29 -342
rect 132 -347 136 -343
rect 42 -363 46 -359
rect 58 -363 62 -359
rect 74 -363 78 -359
rect 90 -363 94 -359
rect 106 -363 110 -359
rect 122 -363 126 -359
rect 132 -377 136 -373
rect 34 -388 38 -384
rect 50 -388 54 -384
rect 66 -388 70 -384
rect 82 -388 86 -384
rect 98 -388 102 -384
rect 114 -388 118 -384
rect 151 -183 155 -179
rect 179 -183 183 -179
rect 193 -183 197 -179
rect 224 -191 228 -187
rect 444 6 448 10
rect 455 -5 459 -1
rect 455 -13 459 -9
rect 455 -21 459 -17
rect 455 -29 459 -25
rect 455 -37 459 -33
rect 455 -45 459 -41
rect 455 -53 459 -49
rect 455 -61 459 -57
rect 455 -69 459 -65
rect 455 -77 459 -73
rect 449 -98 453 -94
rect 455 -116 459 -112
rect 455 -124 459 -120
rect 455 -132 459 -128
rect 455 -140 459 -136
rect 455 -148 459 -144
rect 455 -156 459 -152
rect 455 -164 459 -160
rect 546 6 550 10
rect 558 -5 562 -1
rect 558 -13 562 -9
rect 558 -21 562 -17
rect 558 -29 562 -25
rect 558 -37 562 -33
rect 558 -45 562 -41
rect 558 -53 562 -49
rect 558 -61 562 -57
rect 558 -69 562 -65
rect 558 -77 562 -73
rect 551 -98 555 -94
rect 558 -116 562 -112
rect 558 -124 562 -120
rect 558 -132 562 -128
rect 558 -140 562 -136
rect 558 -148 562 -144
rect 558 -156 562 -152
rect 558 -164 562 -160
rect 268 -191 272 -187
rect 308 -175 312 -171
rect 347 -173 351 -169
rect 363 -173 367 -169
rect 379 -173 383 -169
rect 395 -173 399 -169
rect 411 -173 415 -169
rect 427 -173 431 -169
rect 465 -173 469 -169
rect 481 -173 485 -169
rect 497 -173 501 -169
rect 513 -173 517 -169
rect 529 -173 533 -169
rect 179 -205 183 -201
rect 315 -183 319 -179
rect 308 -197 312 -193
rect 300 -249 304 -245
rect 158 -315 162 -311
rect 158 -347 162 -343
rect 151 -377 155 -373
rect 308 -368 312 -364
rect 339 -197 343 -193
rect 347 -217 351 -213
rect 363 -217 367 -213
rect 379 -217 383 -213
rect 395 -217 399 -213
rect 411 -217 415 -213
rect 427 -217 431 -213
rect 444 -219 448 -215
rect 465 -217 469 -213
rect 481 -217 485 -213
rect 497 -217 501 -213
rect 513 -217 517 -213
rect 529 -217 533 -213
rect 339 -249 343 -245
rect 355 -285 359 -281
rect 371 -285 375 -281
rect 387 -285 391 -281
rect 403 -285 407 -281
rect 419 -285 423 -281
rect 435 -285 439 -281
rect 473 -285 477 -281
rect 489 -285 493 -281
rect 505 -285 509 -281
rect 521 -285 525 -281
rect 537 -285 541 -281
rect 339 -292 343 -288
rect 347 -347 351 -343
rect 363 -347 367 -343
rect 379 -347 383 -343
rect 395 -347 399 -343
rect 411 -347 415 -343
rect 427 -347 431 -343
rect 444 -347 448 -343
rect 465 -347 469 -343
rect 481 -347 485 -343
rect 497 -347 501 -343
rect 513 -347 517 -343
rect 529 -347 533 -343
rect 339 -368 343 -364
<< metal2 >>
rect 129 23 296 25
rect 9 22 296 23
rect 9 20 133 22
rect 9 12 12 20
rect 9 -88 12 8
rect 9 -175 12 -92
rect 16 -99 20 12
rect 16 -201 20 -103
rect 26 -81 29 1
rect 26 -106 29 -85
rect 34 -88 37 12
rect 42 -88 45 12
rect 50 -88 53 12
rect 58 -88 61 12
rect 66 -88 69 12
rect 74 -88 77 12
rect 82 -88 85 12
rect 90 -88 93 12
rect 98 -88 101 12
rect 106 -88 109 12
rect 114 -88 117 12
rect 122 -88 125 12
rect 293 9 296 22
rect 308 24 338 28
rect 308 19 312 24
rect 334 17 442 20
rect 446 17 548 20
rect 330 9 333 16
rect 293 6 333 9
rect 342 6 444 10
rect 448 6 546 10
rect 156 0 197 3
rect 212 0 231 3
rect 134 -4 148 -3
rect 134 -6 186 -4
rect 145 -7 186 -6
rect 194 -5 197 0
rect 297 -4 333 -1
rect 337 -4 455 -1
rect 459 -4 558 -1
rect 194 -8 231 -5
rect 156 -16 197 -13
rect 265 -13 333 -10
rect 337 -12 455 -9
rect 459 -12 558 -9
rect 212 -16 231 -13
rect 134 -20 148 -19
rect 134 -22 186 -20
rect 145 -23 186 -22
rect 194 -21 197 -16
rect 297 -20 333 -17
rect 337 -20 455 -17
rect 459 -20 558 -17
rect 194 -24 231 -21
rect 156 -32 197 -29
rect 265 -29 333 -26
rect 337 -28 455 -25
rect 459 -28 558 -25
rect 212 -32 231 -29
rect 134 -36 148 -35
rect 134 -38 186 -36
rect 145 -39 186 -38
rect 194 -37 197 -32
rect 297 -36 333 -33
rect 337 -36 455 -33
rect 459 -36 558 -33
rect 194 -40 231 -37
rect 156 -48 197 -45
rect 265 -45 333 -42
rect 337 -44 455 -41
rect 459 -44 558 -41
rect 212 -48 231 -45
rect 134 -52 148 -51
rect 134 -54 186 -52
rect 145 -55 186 -54
rect 194 -53 197 -48
rect 297 -52 333 -49
rect 337 -52 455 -49
rect 459 -52 558 -49
rect 194 -56 231 -53
rect 156 -64 197 -61
rect 265 -61 333 -58
rect 337 -60 455 -57
rect 459 -60 558 -57
rect 212 -64 231 -61
rect 134 -68 148 -67
rect 134 -70 186 -68
rect 145 -71 186 -70
rect 194 -69 197 -64
rect 297 -68 333 -65
rect 337 -68 455 -65
rect 459 -68 558 -65
rect 194 -72 231 -69
rect 265 -77 333 -74
rect 337 -76 455 -73
rect 459 -76 558 -73
rect 26 -168 29 -110
rect 34 -173 37 -92
rect 42 -173 45 -92
rect 50 -173 53 -92
rect 58 -173 61 -92
rect 66 -173 69 -92
rect 74 -173 77 -92
rect 82 -173 85 -92
rect 90 -173 93 -92
rect 98 -173 101 -92
rect 106 -173 109 -92
rect 114 -173 117 -92
rect 122 -173 125 -92
rect 319 -98 449 -94
rect 453 -98 551 -94
rect 156 -111 197 -108
rect 212 -111 231 -108
rect 134 -115 148 -114
rect 134 -117 186 -115
rect 145 -118 186 -117
rect 194 -116 197 -111
rect 297 -115 333 -112
rect 337 -115 455 -112
rect 459 -115 558 -112
rect 194 -119 231 -116
rect 156 -127 197 -124
rect 265 -124 333 -121
rect 337 -123 455 -120
rect 459 -123 558 -120
rect 212 -127 231 -124
rect 134 -131 148 -130
rect 134 -133 186 -131
rect 145 -134 186 -133
rect 194 -132 197 -127
rect 297 -131 333 -128
rect 337 -131 455 -128
rect 459 -131 558 -128
rect 194 -135 231 -132
rect 156 -143 197 -140
rect 265 -140 333 -137
rect 337 -139 455 -136
rect 459 -139 558 -136
rect 212 -143 231 -140
rect 134 -147 148 -146
rect 134 -149 186 -147
rect 145 -150 186 -149
rect 194 -148 197 -143
rect 297 -147 333 -144
rect 337 -147 455 -144
rect 459 -147 558 -144
rect 194 -151 231 -148
rect 265 -156 333 -153
rect 337 -155 455 -152
rect 459 -155 558 -152
rect 212 -159 231 -156
rect 134 -163 148 -162
rect 134 -165 186 -163
rect 145 -166 186 -165
rect 297 -163 333 -160
rect 337 -163 455 -160
rect 459 -163 558 -160
rect 34 -176 38 -173
rect 42 -176 46 -173
rect 50 -176 54 -173
rect 58 -176 62 -173
rect 66 -176 70 -173
rect 74 -176 78 -173
rect 82 -176 86 -173
rect 90 -176 94 -173
rect 98 -176 102 -173
rect 106 -176 110 -173
rect 114 -176 118 -173
rect 122 -176 126 -173
rect 173 -175 308 -172
rect 35 -180 38 -176
rect 43 -180 46 -176
rect 51 -180 54 -176
rect 59 -180 62 -176
rect 67 -180 70 -176
rect 75 -180 78 -176
rect 83 -180 86 -176
rect 91 -180 94 -176
rect 99 -180 102 -176
rect 107 -180 110 -176
rect 115 -180 118 -176
rect 123 -180 126 -176
rect 136 -183 151 -180
rect 183 -183 193 -179
rect 197 -183 315 -179
rect 35 -225 38 -184
rect 43 -261 46 -184
rect 51 -225 54 -184
rect 59 -261 62 -184
rect 67 -225 70 -184
rect 75 -261 78 -184
rect 83 -225 86 -184
rect 91 -261 94 -184
rect 99 -225 102 -184
rect 107 -261 110 -184
rect 115 -225 118 -184
rect 123 -261 126 -184
rect 147 -191 224 -187
rect 228 -191 268 -187
rect 312 -197 339 -194
rect 136 -205 179 -201
rect 347 -206 350 -173
rect 363 -206 366 -173
rect 379 -206 382 -173
rect 395 -206 398 -173
rect 411 -206 414 -173
rect 427 -206 430 -173
rect 465 -206 468 -173
rect 481 -206 484 -173
rect 497 -206 500 -173
rect 513 -206 516 -173
rect 529 -206 532 -173
rect 347 -209 359 -206
rect 363 -209 375 -206
rect 379 -209 391 -206
rect 395 -209 407 -206
rect 411 -209 423 -206
rect 427 -209 439 -206
rect 465 -209 477 -206
rect 481 -209 493 -206
rect 497 -209 509 -206
rect 513 -209 525 -206
rect 529 -209 541 -206
rect 304 -249 339 -246
rect 43 -283 46 -265
rect 59 -283 62 -265
rect 75 -283 78 -265
rect 91 -283 94 -265
rect 107 -283 110 -265
rect 123 -283 126 -265
rect 34 -286 46 -283
rect 50 -286 62 -283
rect 66 -286 78 -283
rect 82 -286 94 -283
rect 98 -286 110 -283
rect 114 -286 126 -283
rect 5 -292 25 -288
rect 34 -300 37 -286
rect 50 -300 53 -286
rect 66 -300 69 -286
rect 82 -300 85 -286
rect 98 -300 101 -286
rect 114 -300 117 -286
rect 147 -292 339 -288
rect 41 -308 44 -304
rect 57 -308 60 -304
rect 73 -308 76 -304
rect 89 -308 92 -304
rect 105 -308 108 -304
rect 121 -308 124 -304
rect 12 -314 25 -311
rect 34 -311 44 -308
rect 50 -311 60 -308
rect 66 -311 76 -308
rect 82 -311 92 -308
rect 98 -311 108 -308
rect 114 -311 124 -308
rect 5 -322 25 -318
rect 34 -332 37 -311
rect 12 -346 25 -343
rect 34 -384 37 -336
rect 42 -359 45 -329
rect 50 -332 53 -311
rect 42 -387 45 -363
rect 50 -384 53 -336
rect 58 -359 61 -329
rect 66 -332 69 -311
rect 58 -387 61 -363
rect 66 -384 69 -336
rect 74 -359 77 -329
rect 82 -332 85 -311
rect 74 -387 77 -363
rect 82 -384 85 -336
rect 90 -359 93 -329
rect 98 -332 101 -311
rect 90 -399 93 -363
rect 98 -384 101 -336
rect 106 -359 109 -329
rect 114 -332 117 -311
rect 136 -315 158 -312
rect 347 -316 350 -217
rect 356 -281 359 -209
rect 363 -316 366 -217
rect 372 -281 375 -209
rect 379 -316 382 -217
rect 388 -281 391 -209
rect 395 -316 398 -217
rect 404 -281 407 -209
rect 411 -316 414 -217
rect 420 -281 423 -209
rect 427 -316 430 -217
rect 436 -281 439 -209
rect 347 -319 358 -316
rect 363 -319 374 -316
rect 379 -319 390 -316
rect 395 -319 406 -316
rect 411 -319 422 -316
rect 427 -319 438 -316
rect 106 -393 109 -363
rect 114 -384 117 -336
rect 122 -359 125 -329
rect 136 -347 158 -344
rect 122 -387 125 -363
rect 312 -367 339 -364
rect 136 -376 151 -373
rect 347 -387 350 -347
rect 122 -390 350 -387
rect 355 -393 358 -319
rect 106 -396 358 -393
rect 363 -399 366 -347
rect 371 -384 374 -319
rect 379 -384 382 -347
rect 387 -384 390 -319
rect 395 -384 398 -347
rect 403 -384 406 -319
rect 411 -384 414 -347
rect 419 -384 422 -319
rect 427 -384 430 -347
rect 435 -384 438 -319
rect 444 -343 448 -219
rect 465 -316 468 -217
rect 474 -281 477 -209
rect 481 -316 484 -217
rect 490 -281 493 -209
rect 497 -316 500 -217
rect 506 -281 509 -209
rect 513 -316 516 -217
rect 522 -281 525 -209
rect 529 -316 532 -217
rect 538 -281 541 -209
rect 465 -319 476 -316
rect 481 -319 492 -316
rect 497 -319 508 -316
rect 513 -319 524 -316
rect 529 -319 540 -316
rect 465 -384 468 -347
rect 473 -384 476 -319
rect 481 -384 484 -347
rect 489 -384 492 -319
rect 497 -384 500 -347
rect 505 -384 508 -319
rect 513 -384 516 -347
rect 521 -384 524 -319
rect 529 -384 532 -347
rect 537 -384 540 -319
rect 90 -402 366 -399
<< labels >>
rlabel metal2 42 -365 45 -365 1 RESET
rlabel metal2 58 -365 61 -365 1 load
rlabel metal2 74 -365 77 -365 1 iter
rlabel metal2 90 -365 93 -365 1 InSt0*
rlabel metal2 106 -365 109 -365 1 InSt1*
rlabel metal2 122 -365 125 -365 1 InSt2*
rlabel metal1 300 -383 303 -383 1 p1-
rlabel metal1 308 -383 311 -383 1 p1
rlabel metal1 159 -386 162 -386 1 p2-
rlabel metal1 151 -386 154 -386 1 p2
rlabel metal1 139 -386 147 -386 1 Vdd!
rlabel metal1 315 -383 323 -383 1 GND!
rlabel metal1 347 -341 350 -341 1 OutSt2*
rlabel metal2 355 -341 358 -341 1 OutSt1*
rlabel metal1 363 -341 366 -341 1 OutSt0*
rlabel metal2 371 -341 374 -341 1 ready
rlabel metal1 379 -341 382 -341 1 xr0
rlabel metal2 387 -341 390 -341 1 xr1
rlabel metal1 395 -341 398 -341 1 xw
rlabel metal2 403 -341 406 -341 1 yr0
rlabel metal1 411 -341 414 -341 1 yr1
rlabel metal2 419 -341 422 -341 1 yw
rlabel metal1 427 -341 430 -341 1 osu
rlabel metal2 435 -341 438 -341 1 oss
rlabel metal1 465 -341 468 -341 1 ros
rlabel metal2 473 -341 476 -341 1 g0
rlabel metal1 481 -341 484 -341 1 g1
rlabel metal2 489 -341 492 -341 1 g2
rlabel metal1 497 -341 500 -341 1 g3
rlabel metal2 505 -341 508 -341 1 rfb
rlabel metal1 513 -341 516 -341 1 cin
rlabel metal2 521 -341 524 -341 1 ras
rlabel metal1 529 -341 532 -341 1 ld
rlabel metal2 537 -341 540 -341 1 rd
<< end >>
