magic
tech scmos
timestamp 1003868786
<< error_p >>
rect 156 487 158 507
rect 163 503 164 507
rect 163 487 164 491
rect 196 490 197 494
rect 219 490 221 502
rect 227 490 228 494
rect 84 480 85 484
rect 89 476 91 484
rect 120 480 121 484
rect 84 464 85 468
rect 101 464 103 476
rect 192 467 193 471
rect 231 467 232 471
rect 278 396 282 397
rect 302 396 306 397
rect 326 396 330 397
rect 350 396 354 397
rect 25 381 29 382
rect 57 381 61 382
rect 286 378 298 380
rect 334 378 346 380
rect 25 377 29 378
rect 57 377 61 378
rect 1 367 6 369
rect 17 367 29 369
rect 33 367 37 369
rect 49 367 61 369
rect 65 367 69 369
rect 25 342 29 343
rect 57 342 61 343
rect 25 338 29 339
rect 57 338 61 339
rect 278 338 282 339
rect 302 338 306 339
rect 326 338 330 339
rect 350 338 354 339
rect 504 336 505 338
rect 508 337 509 340
rect 508 336 512 337
rect 520 336 521 338
rect 524 337 525 340
rect 524 336 528 337
rect 536 336 537 338
rect 540 337 541 340
rect 540 336 544 337
rect 584 336 585 338
rect 588 337 589 340
rect 588 336 592 337
rect 600 336 601 338
rect 604 337 605 340
rect 604 336 608 337
rect 616 336 617 338
rect 620 337 621 340
rect 620 336 624 337
rect 632 336 633 338
rect 636 337 637 340
rect 636 336 640 337
rect 648 336 649 338
rect 652 337 653 340
rect 652 336 656 337
rect 504 332 505 333
rect 520 332 521 333
rect 536 332 537 333
rect 584 332 585 333
rect 600 332 601 333
rect 616 332 617 333
rect 632 332 633 333
rect 648 332 649 333
rect 506 326 507 330
rect 522 326 523 330
rect 538 326 539 330
rect 554 326 555 330
rect 570 326 571 330
rect 586 326 587 330
rect 602 326 603 330
rect 618 326 619 330
rect 634 326 635 330
rect 650 326 651 330
rect 666 326 667 330
rect 26 318 27 322
rect 30 319 31 323
rect 58 318 59 322
rect 62 319 63 323
rect 56 305 60 306
rect 492 304 496 305
rect 520 304 521 306
rect 524 305 525 308
rect 524 304 528 305
rect 536 304 537 306
rect 540 305 541 308
rect 540 304 544 305
rect 552 304 553 306
rect 556 305 557 308
rect 556 304 560 305
rect 568 304 569 306
rect 572 305 573 308
rect 572 304 576 305
rect 584 304 585 306
rect 588 305 589 308
rect 588 304 592 305
rect 600 304 601 306
rect 604 305 605 308
rect 604 304 608 305
rect 616 304 617 306
rect 620 305 621 308
rect 620 304 624 305
rect 632 304 633 306
rect 636 305 637 308
rect 636 304 640 305
rect 648 304 649 306
rect 652 305 653 308
rect 652 304 656 305
rect 520 300 521 301
rect 536 300 537 301
rect 552 300 553 301
rect 568 300 569 301
rect 584 300 585 301
rect 600 300 601 301
rect 616 300 617 301
rect 632 300 633 301
rect 648 300 649 301
rect 38 297 39 299
rect 70 297 71 299
rect 31 295 39 297
rect 63 295 71 297
rect 262 296 274 298
rect 310 296 322 298
rect 506 294 507 298
rect 522 294 523 298
rect 538 294 539 298
rect 554 294 555 298
rect 570 294 571 298
rect 586 294 587 298
rect 602 294 603 298
rect 618 294 619 298
rect 634 294 635 298
rect 650 294 651 298
rect 666 294 667 298
rect 38 281 39 285
rect 70 281 71 285
rect 60 278 63 279
rect 506 278 507 282
rect 522 278 523 282
rect 538 278 539 282
rect 554 278 555 282
rect 570 278 571 282
rect 586 278 587 282
rect 602 278 603 282
rect 618 278 619 282
rect 634 278 635 282
rect 650 278 651 282
rect 666 278 667 282
rect 520 275 521 276
rect 536 275 537 276
rect 552 275 553 276
rect 568 275 569 276
rect 584 275 585 276
rect 600 275 601 276
rect 616 275 617 276
rect 632 275 633 276
rect 648 275 649 276
rect 56 274 60 275
rect 492 271 496 272
rect 520 270 521 272
rect 524 271 528 272
rect 278 268 282 269
rect 326 268 330 269
rect 524 268 525 271
rect 536 270 537 272
rect 540 271 544 272
rect 540 268 541 271
rect 552 270 553 272
rect 556 271 560 272
rect 556 268 557 271
rect 568 270 569 272
rect 572 271 576 272
rect 572 268 573 271
rect 584 270 585 272
rect 588 271 592 272
rect 588 268 589 271
rect 600 270 601 272
rect 604 271 608 272
rect 604 268 605 271
rect 616 270 617 272
rect 620 271 624 272
rect 620 268 621 271
rect 632 270 633 272
rect 636 271 640 272
rect 636 268 637 271
rect 648 270 649 272
rect 652 271 656 272
rect 652 268 653 271
<< ntransistor >>
rect 739 718 743 720
rect 840 713 850 715
rect 731 710 735 712
rect 885 652 889 654
rect 901 644 905 646
rect 909 644 913 646
rect 699 636 703 638
rect 710 628 714 630
rect 860 623 870 625
rect 444 578 446 582
rect 444 570 446 574
rect 444 562 446 566
rect 444 554 446 558
rect 444 546 446 550
rect 444 538 446 542
rect 476 578 478 582
rect 476 570 478 574
rect 484 554 486 558
rect 500 570 502 574
rect 492 546 494 550
rect 516 578 518 582
rect 540 578 542 582
rect 540 570 542 574
rect 532 538 534 542
rect 548 562 550 566
rect 612 578 614 582
rect 604 570 606 574
rect 596 562 598 566
rect 596 554 598 558
rect 596 546 598 550
rect 596 538 598 542
rect 628 562 630 566
rect 628 554 630 558
rect 628 546 630 550
rect 620 538 622 542
rect 644 562 646 566
rect 652 562 654 566
rect 644 554 646 558
rect 652 554 654 558
rect 644 546 646 550
rect 652 546 654 550
rect 644 538 646 542
rect 939 620 943 622
rect 947 620 951 622
rect 939 581 943 583
rect 947 581 951 583
rect 939 573 943 575
rect 947 573 951 575
rect 699 557 703 559
rect 885 565 889 567
rect 860 560 870 562
rect 739 557 743 559
rect 710 549 714 551
rect 885 557 889 559
rect 840 552 850 554
rect 731 549 735 551
rect 660 538 662 542
rect 885 549 889 551
rect 860 544 870 546
rect 901 541 905 543
rect 909 541 913 543
rect 16 506 18 510
rect 24 506 26 510
rect 16 498 18 502
rect 24 498 26 502
rect 16 490 18 494
rect 24 490 26 494
rect 16 482 18 486
rect 24 482 26 486
rect 16 474 18 478
rect 24 474 26 478
rect 16 466 18 470
rect 16 458 18 462
rect 48 498 50 502
rect 48 490 50 494
rect 48 482 50 486
rect 48 474 50 478
rect 32 466 34 470
rect 40 466 42 470
rect 64 506 66 510
rect 56 466 58 470
rect 48 458 50 462
rect 56 458 58 462
rect 134 500 138 502
rect 219 495 224 497
rect 142 492 146 494
rect 444 499 446 503
rect 444 491 446 495
rect 444 483 446 487
rect 113 477 117 479
rect 588 491 590 495
rect 596 483 598 487
rect 628 499 630 503
rect 636 499 638 503
rect 628 491 630 495
rect 628 483 630 487
rect 644 483 646 487
rect 699 510 703 512
rect 739 510 743 512
rect 660 499 662 503
rect 710 502 714 504
rect 840 505 850 507
rect 731 502 735 504
rect 660 491 662 495
rect 885 502 889 504
rect 860 497 870 499
rect 739 494 743 496
rect 660 483 662 487
rect 885 494 889 496
rect 840 489 850 491
rect 731 486 735 488
rect 893 486 897 488
rect 955 486 959 488
rect 101 469 105 471
rect 234 464 239 466
rect 8 419 10 423
rect 16 419 18 423
rect 8 411 10 415
rect 64 419 66 423
rect 254 422 258 424
rect 310 422 314 424
rect 350 422 354 424
rect 358 422 362 424
rect 64 411 66 415
rect 254 414 258 416
rect 270 414 274 416
rect 278 414 282 416
rect 286 414 290 416
rect 294 414 298 416
rect 302 414 306 416
rect 310 414 314 416
rect 318 414 322 416
rect 326 414 330 416
rect 334 414 338 416
rect 342 414 346 416
rect 358 414 362 416
rect 30 384 32 391
rect 22 367 24 374
rect 62 384 64 391
rect 299 387 301 393
rect 347 387 349 393
rect 466 450 468 463
rect 458 427 460 440
rect 54 367 56 374
rect 291 378 293 384
rect 498 450 500 463
rect 490 427 492 440
rect 514 450 516 463
rect 506 427 508 440
rect 530 450 532 463
rect 522 427 524 440
rect 546 450 548 463
rect 538 427 540 440
rect 562 450 564 463
rect 554 427 556 440
rect 578 450 580 463
rect 570 427 572 440
rect 594 450 596 463
rect 586 427 588 440
rect 610 450 612 463
rect 602 427 604 440
rect 626 450 628 463
rect 618 427 620 440
rect 642 450 644 463
rect 634 427 636 440
rect 658 450 660 463
rect 952 453 954 465
rect 1038 453 1040 465
rect 650 427 652 440
rect 944 440 946 450
rect 1077 450 1079 463
rect 1069 428 1071 440
rect 267 280 269 286
rect 31 278 35 280
rect 63 278 67 280
rect 890 286 892 298
rect 63 270 67 272
rect 275 271 277 277
rect 323 271 325 277
rect 467 275 471 277
rect 499 275 503 277
rect 515 275 519 277
rect 531 275 535 277
rect 547 275 551 277
rect 563 275 567 277
rect 579 275 583 277
rect 595 275 599 277
rect 611 275 615 277
rect 627 275 631 277
rect 643 275 647 277
rect 659 275 663 277
rect 467 270 471 272
rect 499 270 503 272
rect 515 270 519 272
rect 531 270 535 272
rect 547 270 551 272
rect 563 270 567 272
rect 579 270 583 272
rect 595 270 599 272
rect 611 270 615 272
rect 627 270 631 272
rect 643 270 647 272
rect 659 270 663 272
rect 898 271 900 283
rect 1008 271 1010 283
rect 1078 278 1082 280
<< ptransistor >>
rect 755 718 759 720
rect 808 713 828 715
rect 755 710 759 712
rect 885 684 889 686
rect 893 684 897 686
rect 901 684 905 686
rect 909 684 913 686
rect 939 684 943 686
rect 947 684 951 686
rect 955 684 959 686
rect 683 636 687 638
rect 683 628 687 630
rect 778 623 798 625
rect 254 533 258 535
rect 262 533 266 535
rect 270 533 274 535
rect 278 533 282 535
rect 296 533 300 535
rect 304 533 308 535
rect 360 533 364 535
rect 368 533 372 535
rect 420 578 422 582
rect 420 570 422 574
rect 420 562 422 566
rect 420 554 422 558
rect 420 546 422 550
rect 420 538 422 542
rect 683 557 687 559
rect 778 560 798 562
rect 755 557 759 559
rect 683 549 687 551
rect 808 552 828 554
rect 755 549 759 551
rect 778 544 798 546
rect -16 506 -14 510
rect -16 498 -14 502
rect -16 490 -14 494
rect -16 482 -14 486
rect -16 474 -14 478
rect -16 466 -14 470
rect -16 458 -14 462
rect 156 500 160 502
rect 199 495 209 497
rect 156 492 160 494
rect 87 477 91 479
rect 420 499 422 503
rect 420 491 422 495
rect 420 483 422 487
rect 683 510 687 512
rect 755 510 759 512
rect 683 502 687 504
rect 808 505 828 507
rect 755 502 759 504
rect 778 497 798 499
rect 755 494 759 496
rect 808 489 828 491
rect 755 486 759 488
rect 87 469 91 471
rect 179 464 189 466
rect -16 419 -14 423
rect -16 411 -14 415
rect 22 345 24 357
rect 458 390 460 415
rect 54 345 56 357
rect 30 323 32 335
rect 291 356 293 368
rect 62 323 64 335
rect 490 390 492 415
rect 466 354 468 380
rect 506 390 508 415
rect 498 354 500 380
rect 522 390 524 415
rect 514 354 516 380
rect 538 390 540 415
rect 530 354 532 380
rect 554 390 556 415
rect 546 354 548 380
rect 570 390 572 415
rect 562 354 564 380
rect 586 390 588 415
rect 578 354 580 380
rect 602 390 604 415
rect 594 354 596 380
rect 618 390 620 415
rect 610 354 612 380
rect 634 390 636 415
rect 626 354 628 380
rect 650 390 652 415
rect 642 354 644 380
rect 944 404 946 428
rect 658 354 660 380
rect 299 341 301 353
rect 347 341 349 353
rect 467 336 471 338
rect 499 336 503 338
rect 515 336 519 338
rect 531 336 535 338
rect 547 336 551 338
rect 563 336 567 338
rect 579 336 583 338
rect 595 336 599 338
rect 611 336 615 338
rect 627 336 631 338
rect 643 336 647 338
rect 659 336 663 338
rect 467 331 471 333
rect 499 331 503 333
rect 515 331 519 333
rect 531 331 535 333
rect 547 331 551 333
rect 563 331 567 333
rect 579 331 583 333
rect 595 331 599 333
rect 611 331 615 333
rect 627 331 631 333
rect 643 331 647 333
rect 659 331 663 333
rect 952 377 954 401
rect 1038 377 1040 401
rect 1069 390 1071 416
rect 898 336 900 360
rect 1008 336 1010 360
rect 1077 354 1079 380
rect 275 312 277 324
rect 323 312 325 324
rect 63 305 67 307
rect 31 300 35 302
rect 63 300 67 302
rect 267 296 269 308
rect 467 304 471 306
rect 499 304 503 306
rect 515 304 519 306
rect 531 304 535 306
rect 547 304 551 306
rect 563 304 567 306
rect 579 304 583 306
rect 595 304 599 306
rect 611 304 615 306
rect 627 304 631 306
rect 643 304 647 306
rect 890 310 892 332
rect 659 304 663 306
rect 467 299 471 301
rect 499 299 503 301
rect 515 299 519 301
rect 531 299 535 301
rect 547 299 551 301
rect 563 299 567 301
rect 579 299 583 301
rect 595 299 599 301
rect 611 299 615 301
rect 627 299 631 301
rect 643 299 647 301
rect 659 299 663 301
rect 1078 331 1082 333
rect 1078 302 1082 304
<< ndiffusion >>
rect 739 720 743 721
rect 739 716 743 718
rect 731 713 743 716
rect 731 712 735 713
rect 840 715 850 716
rect 731 709 735 710
rect 840 712 850 713
rect 852 708 853 712
rect 881 655 918 659
rect 935 655 964 659
rect 885 654 889 655
rect 885 651 889 652
rect 901 646 905 647
rect 909 646 913 647
rect 901 643 905 644
rect 909 643 913 644
rect 881 639 918 643
rect 935 639 964 643
rect 699 638 703 639
rect 699 634 703 636
rect 699 631 714 634
rect 710 630 714 631
rect 710 627 714 628
rect 710 624 713 627
rect 852 626 853 630
rect 857 626 858 630
rect 868 626 870 630
rect 860 625 870 626
rect 881 623 918 627
rect 935 623 964 627
rect 860 622 870 623
rect 939 622 943 623
rect 947 622 951 623
rect 447 582 451 585
rect 443 578 444 582
rect 446 578 451 582
rect 447 574 451 578
rect 443 570 444 574
rect 446 570 451 574
rect 447 566 451 570
rect 443 562 444 566
rect 446 562 451 566
rect 447 558 451 562
rect 443 554 444 558
rect 446 554 451 558
rect 447 550 451 554
rect 443 546 444 550
rect 446 546 451 550
rect 447 542 451 546
rect 443 538 444 542
rect 446 538 451 542
rect 447 535 451 538
rect 463 535 467 585
rect 479 582 483 585
rect 475 578 476 582
rect 478 578 483 582
rect 479 574 483 578
rect 475 570 476 574
rect 478 570 483 574
rect 479 558 483 570
rect 479 554 484 558
rect 486 554 487 558
rect 479 535 483 554
rect 495 574 499 585
rect 495 570 500 574
rect 502 570 503 574
rect 495 550 499 570
rect 491 546 492 550
rect 494 546 499 550
rect 495 535 499 546
rect 511 582 515 585
rect 511 578 516 582
rect 518 578 519 582
rect 511 535 515 578
rect 527 542 531 585
rect 543 582 547 585
rect 539 578 540 582
rect 542 578 547 582
rect 543 574 547 578
rect 539 570 540 574
rect 542 570 547 574
rect 527 538 532 542
rect 534 538 535 542
rect 527 535 531 538
rect 543 566 547 570
rect 543 562 548 566
rect 550 562 551 566
rect 543 535 547 562
rect 559 535 563 585
rect 575 535 579 585
rect 591 566 595 585
rect 607 582 611 585
rect 607 578 612 582
rect 614 578 615 582
rect 607 574 611 578
rect 603 570 604 574
rect 606 570 611 574
rect 591 562 596 566
rect 598 562 599 566
rect 591 558 595 562
rect 591 554 596 558
rect 598 554 599 558
rect 591 550 595 554
rect 591 546 596 550
rect 598 546 599 550
rect 591 542 595 546
rect 591 538 596 542
rect 598 538 599 542
rect 591 535 595 538
rect 607 535 611 570
rect 623 566 627 585
rect 623 562 628 566
rect 630 562 631 566
rect 623 558 627 562
rect 623 554 628 558
rect 630 554 631 558
rect 623 550 627 554
rect 623 546 628 550
rect 630 546 631 550
rect 623 542 627 546
rect 619 538 620 542
rect 622 538 627 542
rect 623 535 627 538
rect 639 566 643 585
rect 655 566 659 585
rect 639 562 644 566
rect 646 562 647 566
rect 651 562 652 566
rect 654 562 659 566
rect 639 558 643 562
rect 655 558 659 562
rect 639 554 644 558
rect 646 554 647 558
rect 651 554 652 558
rect 654 554 659 558
rect 639 550 643 554
rect 655 550 659 554
rect 639 546 644 550
rect 646 546 647 550
rect 651 546 652 550
rect 654 546 659 550
rect 639 542 643 546
rect 639 538 644 542
rect 646 538 647 542
rect 639 535 643 538
rect 655 542 659 546
rect 939 619 943 620
rect 947 619 951 620
rect 939 583 943 584
rect 947 583 951 584
rect 881 576 918 580
rect 939 580 943 581
rect 947 580 951 581
rect 935 576 964 580
rect 939 575 943 576
rect 947 575 951 576
rect 939 572 943 573
rect 947 572 951 573
rect 710 561 713 564
rect 699 559 703 560
rect 699 555 703 557
rect 739 559 743 560
rect 840 567 850 568
rect 885 567 889 568
rect 852 563 853 567
rect 857 563 858 567
rect 868 563 870 567
rect 885 564 889 565
rect 860 562 870 563
rect 881 560 918 564
rect 935 560 964 564
rect 996 562 1001 566
rect 860 559 870 560
rect 885 559 889 560
rect 739 555 743 557
rect 699 552 714 555
rect 710 551 714 552
rect 731 552 743 555
rect 731 551 735 552
rect 885 556 889 557
rect 840 554 850 555
rect 655 538 660 542
rect 662 538 663 542
rect 710 548 714 549
rect 731 548 735 549
rect 710 545 713 548
rect 840 551 850 552
rect 885 551 889 552
rect 852 547 853 551
rect 857 547 858 551
rect 868 547 870 551
rect 885 548 889 549
rect 860 546 870 547
rect 881 544 918 548
rect 935 544 964 548
rect 996 546 1001 550
rect 860 543 870 544
rect 901 543 905 544
rect 909 543 913 544
rect 901 540 905 541
rect 655 535 659 538
rect 909 540 913 541
rect 11 510 15 513
rect 27 510 31 513
rect 11 506 16 510
rect 18 506 19 510
rect 23 506 24 510
rect 26 506 31 510
rect 11 502 15 506
rect 27 502 31 506
rect 11 498 16 502
rect 18 498 19 502
rect 23 498 24 502
rect 26 498 31 502
rect 11 494 15 498
rect 27 494 31 498
rect 11 490 16 494
rect 18 490 19 494
rect 23 490 24 494
rect 26 490 31 494
rect 11 486 15 490
rect 27 486 31 490
rect 11 482 16 486
rect 18 482 19 486
rect 23 482 24 486
rect 26 482 31 486
rect 11 478 15 482
rect 27 478 31 482
rect 11 474 16 478
rect 18 474 19 478
rect 23 474 24 478
rect 26 474 31 478
rect 11 470 15 474
rect 11 466 16 470
rect 18 466 19 470
rect 11 462 15 466
rect 11 458 16 462
rect 18 458 19 462
rect 11 455 15 458
rect 27 470 31 474
rect 43 502 47 513
rect 43 498 48 502
rect 50 498 51 502
rect 43 494 47 498
rect 43 490 48 494
rect 50 490 51 494
rect 43 486 47 490
rect 43 482 48 486
rect 50 482 51 486
rect 43 478 47 482
rect 43 474 48 478
rect 50 474 51 478
rect 43 470 47 474
rect 27 466 32 470
rect 34 466 35 470
rect 39 466 40 470
rect 42 466 47 470
rect 27 455 31 466
rect 43 462 47 466
rect 59 510 63 513
rect 59 506 64 510
rect 66 506 67 510
rect 59 470 63 506
rect 55 466 56 470
rect 58 466 63 470
rect 59 462 63 466
rect 43 458 48 462
rect 50 458 51 462
rect 55 458 56 462
rect 58 458 63 462
rect 43 455 47 458
rect 59 455 63 458
rect 134 502 138 503
rect 134 498 138 500
rect 134 495 146 498
rect 142 494 146 495
rect 219 497 224 498
rect 142 491 146 492
rect 219 494 224 495
rect 113 480 116 483
rect 447 503 451 506
rect 443 499 444 503
rect 446 499 451 503
rect 447 495 451 499
rect 443 491 444 495
rect 446 491 451 495
rect 447 487 451 491
rect 443 483 444 487
rect 446 483 451 487
rect 113 479 117 480
rect 113 476 117 477
rect 101 473 117 476
rect 101 471 105 473
rect 447 480 451 483
rect 463 480 467 506
rect 479 480 483 506
rect 495 480 499 506
rect 511 480 515 506
rect 527 480 531 506
rect 543 480 547 506
rect 559 480 563 506
rect 575 480 579 506
rect 591 495 595 506
rect 587 491 588 495
rect 590 491 595 495
rect 591 487 595 491
rect 591 483 596 487
rect 598 483 599 487
rect 591 480 595 483
rect 607 480 611 506
rect 623 503 627 506
rect 639 503 643 506
rect 623 499 628 503
rect 630 499 631 503
rect 635 499 636 503
rect 638 499 643 503
rect 623 495 627 499
rect 623 491 628 495
rect 630 491 631 495
rect 623 487 627 491
rect 623 483 628 487
rect 630 483 631 487
rect 623 480 627 483
rect 639 487 643 499
rect 639 483 644 487
rect 646 483 647 487
rect 639 480 643 483
rect 655 503 659 506
rect 699 512 703 513
rect 699 508 703 510
rect 739 512 743 513
rect 739 508 743 510
rect 699 505 714 508
rect 710 504 714 505
rect 655 499 660 503
rect 662 499 663 503
rect 731 505 743 508
rect 731 504 735 505
rect 840 507 850 508
rect 655 495 659 499
rect 655 491 660 495
rect 662 491 663 495
rect 710 501 714 502
rect 731 501 735 502
rect 710 498 713 501
rect 739 496 743 497
rect 840 504 850 505
rect 885 504 889 505
rect 852 500 853 504
rect 857 500 858 504
rect 868 500 870 504
rect 885 501 889 502
rect 860 499 870 500
rect 881 497 918 501
rect 935 497 964 501
rect 860 496 870 497
rect 885 496 889 497
rect 739 492 743 494
rect 655 487 659 491
rect 655 483 660 487
rect 662 483 663 487
rect 731 489 743 492
rect 731 488 735 489
rect 885 493 889 494
rect 840 491 850 492
rect 731 485 735 486
rect 655 480 659 483
rect 840 488 850 489
rect 893 488 897 489
rect 955 488 959 489
rect 852 484 853 488
rect 893 485 897 486
rect 881 481 918 485
rect 955 485 959 486
rect 935 481 964 485
rect 101 468 105 469
rect 237 467 239 471
rect 234 466 239 467
rect 250 464 367 468
rect 371 464 372 468
rect 901 467 905 468
rect 234 463 239 464
rect 11 423 15 426
rect 7 419 8 423
rect 10 419 16 423
rect 18 419 19 423
rect 11 415 15 419
rect 7 411 8 415
rect 10 411 15 415
rect 11 408 15 411
rect 27 408 31 426
rect 43 408 47 426
rect 59 423 63 426
rect 254 424 258 425
rect 310 424 314 425
rect 350 424 354 425
rect 441 427 442 440
rect 358 424 362 425
rect 59 419 64 423
rect 66 419 67 423
rect 254 421 258 422
rect 310 421 314 422
rect 350 421 354 422
rect 358 421 362 422
rect 59 415 63 419
rect 250 417 367 421
rect 371 417 377 421
rect 254 416 258 417
rect 270 416 274 417
rect 278 416 282 417
rect 286 416 290 417
rect 294 416 298 417
rect 302 416 306 417
rect 310 416 314 417
rect 318 416 322 417
rect 326 416 330 417
rect 334 416 338 417
rect 342 416 346 417
rect 358 416 362 417
rect 59 411 64 415
rect 66 411 67 415
rect 254 413 258 414
rect 59 408 63 411
rect 270 413 274 414
rect 278 413 282 414
rect 286 413 290 414
rect 294 413 298 414
rect 302 413 306 414
rect 310 413 314 414
rect 318 413 322 414
rect 326 413 330 414
rect 334 413 338 414
rect 342 413 346 414
rect 358 413 362 414
rect 25 389 30 391
rect 29 384 30 389
rect 32 384 33 391
rect 57 389 62 391
rect 5 367 6 374
rect 21 367 22 374
rect 24 367 25 374
rect 61 384 62 389
rect 64 384 65 391
rect 278 387 281 392
rect 295 387 299 393
rect 301 392 302 393
rect 301 387 305 392
rect 326 387 329 392
rect 343 387 347 393
rect 349 392 350 393
rect 349 387 353 392
rect 463 461 466 463
rect 465 450 466 461
rect 468 450 469 463
rect 495 461 498 463
rect 461 447 465 448
rect 461 442 465 443
rect 457 427 458 440
rect 460 427 461 440
rect 295 384 298 387
rect 53 367 54 374
rect 56 367 57 374
rect 287 382 291 384
rect 290 378 291 382
rect 293 378 298 384
rect 343 384 346 387
rect 335 382 346 384
rect 338 378 346 382
rect 497 450 498 461
rect 500 450 501 463
rect 511 461 514 463
rect 493 447 497 448
rect 493 442 497 443
rect 489 427 490 440
rect 492 427 493 440
rect 513 450 514 461
rect 516 450 517 463
rect 527 461 530 463
rect 509 447 513 448
rect 509 442 513 443
rect 505 427 506 440
rect 508 427 509 440
rect 529 450 530 461
rect 532 450 533 463
rect 543 461 546 463
rect 525 447 529 448
rect 525 442 529 443
rect 521 427 522 440
rect 524 427 525 440
rect 545 450 546 461
rect 548 450 549 463
rect 559 461 562 463
rect 541 447 545 448
rect 541 442 545 443
rect 537 427 538 440
rect 540 427 541 440
rect 561 450 562 461
rect 564 450 565 463
rect 575 461 578 463
rect 557 447 561 448
rect 557 442 561 443
rect 553 427 554 440
rect 556 427 557 440
rect 577 450 578 461
rect 580 450 581 463
rect 591 461 594 463
rect 573 447 577 448
rect 573 442 577 443
rect 569 427 570 440
rect 572 427 573 440
rect 593 450 594 461
rect 596 450 597 463
rect 607 461 610 463
rect 589 447 593 448
rect 589 442 593 443
rect 585 427 586 440
rect 588 427 589 440
rect 609 450 610 461
rect 612 450 613 463
rect 623 461 626 463
rect 605 447 609 448
rect 605 442 609 443
rect 601 427 602 440
rect 604 427 605 440
rect 625 450 626 461
rect 628 450 629 463
rect 639 461 642 463
rect 621 447 625 448
rect 621 442 625 443
rect 617 427 618 440
rect 620 427 621 440
rect 641 450 642 461
rect 644 450 645 463
rect 655 461 658 463
rect 637 447 641 448
rect 637 442 641 443
rect 633 427 634 440
rect 636 427 637 440
rect 657 450 658 461
rect 660 450 661 463
rect 955 467 959 468
rect 901 453 904 458
rect 948 453 952 465
rect 954 458 955 465
rect 1011 467 1015 468
rect 1074 480 1078 481
rect 1041 467 1045 468
rect 954 453 958 458
rect 1011 453 1014 458
rect 1034 453 1038 465
rect 1040 458 1041 465
rect 1074 461 1077 463
rect 1040 453 1044 458
rect 948 450 951 453
rect 653 447 657 448
rect 653 442 657 443
rect 649 427 650 440
rect 652 427 653 440
rect 940 448 944 450
rect 943 440 944 448
rect 946 440 951 450
rect 1034 450 1037 453
rect 1026 448 1037 450
rect 1029 440 1037 448
rect 1076 450 1077 461
rect 1079 450 1080 463
rect 1072 447 1076 448
rect 1072 442 1076 443
rect 1068 428 1069 440
rect 1071 428 1072 440
rect 31 280 35 281
rect 266 282 267 286
rect 63 280 67 281
rect 263 280 267 282
rect 269 280 274 286
rect 31 277 35 278
rect 63 272 67 278
rect 271 277 274 280
rect 314 282 322 286
rect 311 280 322 282
rect 319 277 322 280
rect 889 288 890 298
rect 886 286 890 288
rect 892 286 897 298
rect 473 278 474 282
rect 467 277 471 278
rect 499 277 503 278
rect 515 277 519 278
rect 531 277 535 278
rect 547 277 551 278
rect 563 277 567 278
rect 579 277 583 278
rect 595 277 599 278
rect 611 277 615 278
rect 627 277 631 278
rect 643 277 647 278
rect 894 283 897 286
rect 999 288 1007 298
rect 956 286 959 288
rect 996 286 1007 288
rect 1004 283 1007 286
rect 1042 286 1045 288
rect 659 277 663 278
rect 271 271 275 277
rect 277 272 281 277
rect 277 271 278 272
rect 63 269 67 270
rect 319 271 323 277
rect 325 272 329 277
rect 467 272 471 275
rect 499 272 503 275
rect 515 272 519 275
rect 531 272 535 275
rect 547 272 551 275
rect 563 272 567 275
rect 579 272 583 275
rect 595 272 599 275
rect 611 272 615 275
rect 627 272 631 275
rect 643 272 647 275
rect 659 272 663 275
rect 325 271 326 272
rect 467 269 471 270
rect 467 266 468 269
rect 499 269 503 270
rect 515 269 519 270
rect 515 267 516 269
rect 531 269 535 270
rect 547 269 551 270
rect 563 269 567 270
rect 579 269 583 270
rect 595 269 599 270
rect 611 269 615 270
rect 627 269 631 270
rect 643 269 647 270
rect 894 271 898 283
rect 900 278 904 283
rect 955 278 958 283
rect 900 271 901 278
rect 659 269 663 270
rect 901 268 905 269
rect 1004 271 1008 283
rect 1010 278 1014 283
rect 1041 278 1044 283
rect 1084 281 1085 285
rect 1078 280 1082 281
rect 1010 271 1011 278
rect 955 268 959 269
rect 1011 268 1015 269
rect 1041 268 1045 269
rect 1078 272 1082 278
<< pdiffusion >>
rect 761 721 762 725
rect 755 720 759 721
rect 755 717 759 718
rect 808 716 813 720
rect 755 712 759 713
rect 808 715 828 716
rect 808 712 828 713
rect 755 709 759 710
rect 761 705 762 709
rect 805 708 806 712
rect 883 691 963 692
rect 885 686 889 687
rect 893 686 897 687
rect 901 686 905 687
rect 909 686 913 687
rect 939 686 943 687
rect 947 686 951 687
rect 955 686 959 687
rect 885 683 889 684
rect 893 683 897 684
rect 901 683 905 684
rect 909 683 913 684
rect 939 683 943 684
rect 947 683 951 684
rect 955 683 959 684
rect 680 639 681 643
rect 683 638 687 639
rect 683 635 687 636
rect 683 630 687 631
rect 683 627 687 628
rect 680 623 681 627
rect 778 626 780 630
rect 800 626 801 630
rect 805 626 806 630
rect 778 625 798 626
rect 778 622 798 623
rect 778 618 780 622
rect 252 540 310 541
rect 254 535 258 536
rect 262 535 266 536
rect 270 535 274 536
rect 278 535 282 536
rect 296 535 300 536
rect 304 535 308 536
rect 360 535 364 536
rect 368 535 372 536
rect 414 536 415 584
rect 419 578 420 582
rect 422 578 423 582
rect 419 570 420 574
rect 422 570 423 574
rect 419 562 420 566
rect 422 562 423 566
rect 419 554 420 558
rect 422 554 423 558
rect 419 546 420 550
rect 422 546 423 550
rect 419 538 420 542
rect 422 538 423 542
rect 254 532 258 533
rect 262 532 266 533
rect 270 532 274 533
rect 278 532 282 533
rect 296 532 300 533
rect 304 532 308 533
rect 360 532 364 533
rect 368 532 372 533
rect 808 567 828 568
rect 680 560 681 564
rect 683 559 687 560
rect 683 556 687 557
rect 761 560 762 564
rect 778 563 780 567
rect 800 563 801 567
rect 805 563 806 567
rect 755 559 759 560
rect 778 562 798 563
rect 778 559 798 560
rect 683 551 687 552
rect 755 556 759 557
rect 778 555 780 559
rect 808 555 813 559
rect 755 551 759 552
rect 808 554 828 555
rect 808 551 828 552
rect 683 548 687 549
rect 680 544 681 548
rect 755 548 759 549
rect 761 544 762 548
rect 778 547 780 551
rect 800 547 801 551
rect 805 547 806 551
rect 778 546 798 547
rect 778 543 798 544
rect 778 539 780 543
rect -22 456 -21 512
rect -17 506 -16 510
rect -14 506 -13 510
rect -17 498 -16 502
rect -14 498 -13 502
rect -17 490 -16 494
rect -14 490 -13 494
rect -17 482 -16 486
rect -14 482 -13 486
rect -17 474 -16 478
rect -14 474 -13 478
rect -17 466 -16 470
rect -14 466 -13 470
rect -17 458 -16 462
rect -14 458 -13 462
rect 156 502 160 503
rect 156 499 160 500
rect 156 494 160 495
rect 199 498 204 502
rect 199 497 209 498
rect 199 494 209 495
rect 156 491 160 492
rect 87 479 91 480
rect 414 481 415 505
rect 419 499 420 503
rect 422 499 423 503
rect 419 491 420 495
rect 422 491 423 495
rect 419 483 420 487
rect 422 483 423 487
rect 87 476 91 477
rect 87 471 91 472
rect 680 513 681 517
rect 683 512 687 513
rect 683 509 687 510
rect 761 513 762 517
rect 755 512 759 513
rect 683 504 687 505
rect 755 509 759 510
rect 808 508 813 512
rect 755 504 759 505
rect 808 507 828 508
rect 808 504 828 505
rect 683 501 687 502
rect 680 497 681 501
rect 755 501 759 502
rect 761 497 762 501
rect 778 500 780 504
rect 800 500 801 504
rect 805 500 806 504
rect 755 496 759 497
rect 778 499 798 500
rect 778 496 798 497
rect 755 493 759 494
rect 778 492 780 496
rect 808 492 813 496
rect 755 488 759 489
rect 808 491 828 492
rect 808 488 828 489
rect 755 485 759 486
rect 761 481 762 485
rect 805 484 806 488
rect 87 468 91 469
rect 179 467 181 471
rect 179 466 189 467
rect 179 463 189 464
rect 179 459 181 463
rect -22 409 -21 425
rect -17 419 -16 423
rect -14 419 -13 423
rect -17 411 -16 415
rect -14 411 -13 415
rect 5 352 6 357
rect 21 352 22 357
rect 3 345 6 352
rect 19 345 22 352
rect 24 345 25 357
rect 441 397 442 415
rect 439 390 442 397
rect 457 397 458 415
rect 455 390 458 397
rect 460 390 461 415
rect 53 352 54 357
rect 51 345 54 352
rect 56 345 57 357
rect 29 325 30 335
rect 25 323 30 325
rect 32 332 33 335
rect 32 323 35 332
rect 290 358 291 368
rect 287 356 291 358
rect 293 356 298 368
rect 61 325 62 335
rect 57 323 62 325
rect 64 332 65 335
rect 64 323 67 332
rect 31 302 35 308
rect 278 348 281 353
rect 295 353 298 356
rect 338 358 346 368
rect 335 356 346 358
rect 343 353 346 356
rect 461 387 465 388
rect 461 382 465 383
rect 489 397 490 415
rect 487 390 490 397
rect 492 390 493 415
rect 465 356 466 380
rect 461 354 466 356
rect 468 363 469 380
rect 468 354 471 363
rect 493 387 497 388
rect 493 382 497 383
rect 505 397 506 415
rect 503 390 506 397
rect 508 390 509 415
rect 497 356 498 380
rect 493 354 498 356
rect 500 363 501 380
rect 500 354 503 363
rect 509 387 513 388
rect 509 382 513 383
rect 521 397 522 415
rect 519 390 522 397
rect 524 390 525 415
rect 513 356 514 380
rect 509 354 514 356
rect 516 363 517 380
rect 516 354 519 363
rect 525 387 529 388
rect 525 382 529 383
rect 537 397 538 415
rect 535 390 538 397
rect 540 390 541 415
rect 529 356 530 380
rect 525 354 530 356
rect 532 363 533 380
rect 532 354 535 363
rect 541 387 545 388
rect 541 382 545 383
rect 553 397 554 415
rect 551 390 554 397
rect 556 390 557 415
rect 545 356 546 380
rect 541 354 546 356
rect 548 363 549 380
rect 548 354 551 363
rect 557 387 561 388
rect 557 382 561 383
rect 569 397 570 415
rect 567 390 570 397
rect 572 390 573 415
rect 561 356 562 380
rect 557 354 562 356
rect 564 363 565 380
rect 564 354 567 363
rect 573 387 577 388
rect 573 382 577 383
rect 585 397 586 415
rect 583 390 586 397
rect 588 390 589 415
rect 577 356 578 380
rect 573 354 578 356
rect 580 363 581 380
rect 580 354 583 363
rect 589 387 593 388
rect 589 382 593 383
rect 601 397 602 415
rect 599 390 602 397
rect 604 390 605 415
rect 593 356 594 380
rect 589 354 594 356
rect 596 363 597 380
rect 596 354 599 363
rect 605 387 609 388
rect 605 382 609 383
rect 617 397 618 415
rect 615 390 618 397
rect 620 390 621 415
rect 609 356 610 380
rect 605 354 610 356
rect 612 363 613 380
rect 612 354 615 363
rect 621 387 625 388
rect 621 382 625 383
rect 633 397 634 415
rect 631 390 634 397
rect 636 390 637 415
rect 625 356 626 380
rect 621 354 626 356
rect 628 363 629 380
rect 628 354 631 363
rect 637 387 641 388
rect 637 382 641 383
rect 649 397 650 415
rect 647 390 650 397
rect 652 390 653 415
rect 641 356 642 380
rect 637 354 642 356
rect 644 363 645 380
rect 644 354 647 363
rect 653 387 657 388
rect 653 382 657 383
rect 943 406 944 428
rect 940 404 944 406
rect 946 404 951 428
rect 657 356 658 380
rect 653 354 658 356
rect 660 363 661 380
rect 660 354 663 363
rect 295 341 299 353
rect 301 348 305 353
rect 326 348 329 353
rect 301 341 302 348
rect 343 341 347 353
rect 349 348 353 353
rect 349 341 350 348
rect 467 339 468 341
rect 467 338 471 339
rect 499 338 503 339
rect 515 338 519 339
rect 531 338 535 339
rect 547 338 551 339
rect 563 339 564 341
rect 563 338 567 339
rect 579 339 580 341
rect 579 338 583 339
rect 595 338 599 339
rect 611 338 615 339
rect 627 338 631 339
rect 643 338 647 339
rect 659 338 663 339
rect 467 333 471 336
rect 499 333 503 336
rect 515 333 519 336
rect 531 333 535 336
rect 547 333 551 336
rect 563 333 567 336
rect 579 333 583 336
rect 595 333 599 336
rect 611 333 615 336
rect 627 333 631 336
rect 643 333 647 336
rect 659 333 663 336
rect 901 396 904 401
rect 948 401 951 404
rect 1029 406 1037 428
rect 1026 404 1037 406
rect 1034 401 1037 404
rect 948 377 952 401
rect 954 396 958 401
rect 1011 396 1014 401
rect 954 377 955 396
rect 901 374 905 375
rect 955 374 959 375
rect 1034 377 1038 401
rect 1040 396 1044 401
rect 1068 397 1069 416
rect 1040 377 1041 396
rect 1066 390 1069 397
rect 1071 390 1072 416
rect 1011 374 1015 375
rect 1041 374 1045 375
rect 894 336 898 360
rect 900 336 901 360
rect 1004 336 1008 360
rect 1010 336 1011 360
rect 1072 387 1076 388
rect 1072 382 1076 383
rect 1076 356 1077 380
rect 1072 354 1077 356
rect 1079 363 1080 380
rect 1079 354 1082 363
rect 894 332 897 336
rect 271 312 275 324
rect 277 312 278 324
rect 319 312 323 324
rect 325 312 326 324
rect 467 330 471 331
rect 473 326 474 330
rect 499 330 503 331
rect 515 330 519 331
rect 531 330 535 331
rect 547 330 551 331
rect 563 330 567 331
rect 579 330 583 331
rect 595 330 599 331
rect 611 330 615 331
rect 627 330 631 331
rect 643 330 647 331
rect 659 330 663 331
rect 271 308 274 312
rect 63 307 67 308
rect 63 302 67 305
rect 31 299 35 300
rect 63 299 67 300
rect 266 296 267 308
rect 269 296 274 308
rect 319 308 322 312
rect 314 296 322 308
rect 467 307 468 309
rect 467 306 471 307
rect 499 306 503 307
rect 515 307 516 309
rect 515 306 519 307
rect 531 306 535 307
rect 547 306 551 307
rect 563 306 567 307
rect 579 306 583 307
rect 595 306 599 307
rect 611 306 615 307
rect 627 306 631 307
rect 643 306 647 307
rect 889 310 890 332
rect 892 310 897 332
rect 659 306 663 307
rect 467 301 471 304
rect 499 301 503 304
rect 515 301 519 304
rect 531 301 535 304
rect 547 301 551 304
rect 563 301 567 304
rect 579 301 583 304
rect 595 301 599 304
rect 611 301 615 304
rect 627 301 631 304
rect 643 301 647 304
rect 659 301 663 304
rect 467 298 471 299
rect 473 294 474 298
rect 499 298 503 299
rect 515 298 519 299
rect 531 298 535 299
rect 547 298 551 299
rect 563 298 567 299
rect 579 298 583 299
rect 595 298 599 299
rect 611 298 615 299
rect 627 298 631 299
rect 643 298 647 299
rect 659 298 663 299
rect 1004 332 1007 336
rect 999 310 1007 332
rect 1078 333 1082 339
rect 1078 330 1082 331
rect 1084 326 1085 330
rect 1078 304 1082 308
rect 1078 301 1082 302
rect 1084 299 1088 301
rect 1084 297 1085 299
<< ndcontact >>
rect 739 721 743 725
rect 840 716 850 720
rect 731 705 735 709
rect 840 708 852 712
rect 901 663 905 667
rect 909 663 913 667
rect 918 655 922 659
rect 964 655 968 659
rect 885 647 889 651
rect 901 647 905 651
rect 909 647 913 651
rect 699 639 703 643
rect 918 639 922 643
rect 964 639 968 643
rect 893 631 897 635
rect 955 631 959 635
rect 713 623 717 627
rect 840 626 852 630
rect 858 626 868 630
rect 918 623 922 627
rect 964 623 968 627
rect 860 618 870 622
rect 447 585 451 589
rect 439 578 443 582
rect 439 570 443 574
rect 439 562 443 566
rect 439 554 443 558
rect 439 546 443 550
rect 439 538 443 542
rect 447 531 451 535
rect 463 585 467 589
rect 463 531 467 535
rect 479 585 483 589
rect 471 578 475 582
rect 471 570 475 574
rect 487 554 491 558
rect 479 531 483 535
rect 495 585 499 589
rect 503 570 507 574
rect 487 546 491 550
rect 495 531 499 535
rect 511 585 515 589
rect 519 578 523 582
rect 511 531 515 535
rect 527 585 531 589
rect 543 585 547 589
rect 535 578 539 582
rect 535 570 539 574
rect 535 538 539 542
rect 527 531 531 535
rect 551 562 555 566
rect 543 531 547 535
rect 559 585 563 589
rect 559 531 563 535
rect 575 585 579 589
rect 575 531 579 535
rect 591 585 595 589
rect 607 585 611 589
rect 615 578 619 582
rect 599 570 603 574
rect 599 562 603 566
rect 599 554 603 558
rect 599 546 603 550
rect 599 538 603 542
rect 591 531 595 535
rect 607 531 611 535
rect 623 585 627 589
rect 631 562 635 566
rect 631 554 635 558
rect 631 546 635 550
rect 615 538 619 542
rect 623 531 627 535
rect 639 585 643 589
rect 655 585 659 589
rect 647 562 651 566
rect 647 554 651 558
rect 647 546 651 550
rect 647 538 651 542
rect 639 531 643 535
rect 939 615 943 619
rect 947 615 951 619
rect 939 584 943 588
rect 947 584 951 588
rect 918 576 922 580
rect 964 576 968 580
rect 885 568 889 572
rect 939 568 943 572
rect 947 568 951 572
rect 699 560 703 564
rect 713 560 717 564
rect 731 560 735 564
rect 739 560 743 564
rect 840 563 852 567
rect 858 563 868 567
rect 918 560 922 564
rect 964 560 968 564
rect 1001 562 1005 566
rect 840 555 850 559
rect 860 555 870 559
rect 885 552 889 556
rect 663 538 667 542
rect 713 544 717 548
rect 731 544 735 548
rect 840 547 852 551
rect 858 547 868 551
rect 918 544 922 548
rect 964 544 968 548
rect 1001 546 1005 550
rect 860 539 870 543
rect 655 531 659 535
rect 901 536 905 540
rect 909 536 913 540
rect 11 513 15 517
rect 27 513 31 517
rect 19 506 23 510
rect 19 498 23 502
rect 19 490 23 494
rect 19 482 23 486
rect 19 474 23 478
rect 19 466 23 470
rect 19 458 23 462
rect 11 451 15 455
rect 43 513 47 517
rect 51 498 55 502
rect 51 490 55 494
rect 51 482 55 486
rect 51 474 55 478
rect 35 466 39 470
rect 27 451 31 455
rect 59 513 63 517
rect 67 506 71 510
rect 51 466 55 470
rect 51 458 55 462
rect 43 451 47 455
rect 59 451 63 455
rect 134 503 138 507
rect 67 489 71 493
rect 219 498 224 502
rect 142 487 146 491
rect 219 490 227 494
rect 116 480 120 484
rect 447 506 451 510
rect 439 499 443 503
rect 439 491 443 495
rect 439 483 443 487
rect 447 476 451 480
rect 463 506 467 510
rect 463 476 467 480
rect 479 506 483 510
rect 479 476 483 480
rect 495 506 499 510
rect 495 476 499 480
rect 511 506 515 510
rect 511 476 515 480
rect 527 506 531 510
rect 527 476 531 480
rect 543 506 547 510
rect 543 476 547 480
rect 559 506 563 510
rect 559 476 563 480
rect 575 506 579 510
rect 575 476 579 480
rect 591 506 595 510
rect 583 491 587 495
rect 599 483 603 487
rect 591 476 595 480
rect 607 506 611 510
rect 607 476 611 480
rect 623 506 627 510
rect 639 506 643 510
rect 631 499 635 503
rect 631 491 635 495
rect 631 483 635 487
rect 623 476 627 480
rect 647 483 651 487
rect 639 476 643 480
rect 655 506 659 510
rect 699 513 703 517
rect 739 513 743 517
rect 663 499 667 503
rect 840 508 850 512
rect 885 505 889 509
rect 663 491 667 495
rect 713 497 717 501
rect 731 497 735 501
rect 739 497 743 501
rect 840 500 852 504
rect 858 500 868 504
rect 918 497 922 501
rect 964 497 968 501
rect 663 483 667 487
rect 840 492 850 496
rect 860 492 870 496
rect 885 489 889 493
rect 893 489 897 493
rect 955 489 959 493
rect 655 476 659 480
rect 731 481 735 485
rect 840 484 852 488
rect 918 481 922 485
rect 964 481 968 485
rect 67 458 71 462
rect 101 464 105 468
rect 231 467 237 471
rect 367 464 371 468
rect 234 459 239 463
rect 11 426 15 430
rect 3 419 7 423
rect 19 419 23 423
rect 3 411 7 415
rect 11 404 15 408
rect 27 426 31 430
rect 27 404 31 408
rect 43 426 47 430
rect 43 404 47 408
rect 59 426 63 430
rect 254 425 258 429
rect 310 425 314 429
rect 350 425 354 429
rect 358 425 362 429
rect 437 427 441 440
rect 67 419 71 423
rect 367 417 371 421
rect 377 417 381 421
rect 67 411 71 415
rect 59 404 63 408
rect 254 409 258 413
rect 270 409 274 413
rect 278 409 282 413
rect 286 409 290 413
rect 294 409 298 413
rect 302 409 306 413
rect 310 409 314 413
rect 318 409 322 413
rect 326 409 330 413
rect 334 409 338 413
rect 342 409 346 413
rect 358 409 362 413
rect 278 392 282 396
rect 25 381 29 389
rect 33 384 37 391
rect 1 367 5 374
rect 17 367 21 374
rect 25 367 29 377
rect 57 381 61 389
rect 65 384 69 391
rect 302 392 306 396
rect 326 392 330 396
rect 350 392 354 396
rect 461 448 465 461
rect 469 450 473 463
rect 485 450 489 463
rect 453 427 457 440
rect 461 427 465 442
rect 33 367 37 374
rect 49 367 53 374
rect 57 367 61 377
rect 286 378 290 382
rect 65 367 69 374
rect 334 378 338 382
rect 493 448 497 461
rect 501 450 505 463
rect 469 427 473 440
rect 485 427 489 440
rect 493 427 497 442
rect 509 448 513 461
rect 517 450 521 463
rect 501 427 505 440
rect 509 427 513 442
rect 525 448 529 461
rect 533 450 537 463
rect 517 427 521 440
rect 525 427 529 442
rect 541 448 545 461
rect 549 450 553 463
rect 533 427 537 440
rect 541 427 545 442
rect 557 448 561 461
rect 565 450 569 463
rect 549 427 553 440
rect 557 427 561 442
rect 573 448 577 461
rect 581 450 585 463
rect 565 427 569 440
rect 573 427 577 442
rect 589 448 593 461
rect 597 450 601 463
rect 581 427 585 440
rect 589 427 593 442
rect 605 448 609 461
rect 613 450 617 463
rect 597 427 601 440
rect 605 427 609 442
rect 621 448 625 461
rect 629 450 633 463
rect 613 427 617 440
rect 621 427 625 442
rect 637 448 641 461
rect 645 450 649 463
rect 629 427 633 440
rect 637 427 641 442
rect 653 448 657 461
rect 661 450 665 463
rect 901 458 905 467
rect 955 458 959 467
rect 1011 458 1015 467
rect 1074 476 1078 480
rect 1041 458 1045 467
rect 645 427 649 440
rect 653 427 657 442
rect 939 440 943 448
rect 661 427 665 440
rect 1025 440 1029 448
rect 1072 448 1076 461
rect 1080 450 1084 463
rect 1064 428 1068 440
rect 1072 428 1076 442
rect 1080 428 1084 440
rect 31 281 38 285
rect 63 281 70 285
rect 262 282 266 286
rect 31 273 35 277
rect 310 282 314 286
rect 885 288 889 298
rect 467 278 473 282
rect 499 278 506 282
rect 515 278 522 282
rect 531 278 538 282
rect 547 278 554 282
rect 563 278 570 282
rect 579 278 586 282
rect 595 278 602 282
rect 611 278 618 282
rect 627 278 634 282
rect 643 278 650 282
rect 659 278 666 282
rect 955 288 959 298
rect 995 288 999 298
rect 1041 288 1045 298
rect 63 265 67 269
rect 278 268 282 272
rect 326 268 330 272
rect 468 265 472 269
rect 499 265 503 269
rect 516 265 520 269
rect 531 265 535 269
rect 547 265 551 269
rect 563 265 567 269
rect 579 265 583 269
rect 595 265 599 269
rect 611 265 615 269
rect 627 265 631 269
rect 643 265 647 269
rect 901 269 905 278
rect 659 265 663 269
rect 955 269 959 278
rect 1078 281 1084 285
rect 1011 269 1015 278
rect 1041 269 1045 278
rect 1078 268 1082 272
<< pdcontact >>
rect 755 721 761 725
rect 755 713 759 717
rect 813 716 828 720
rect 755 705 761 709
rect 806 708 828 712
rect 883 687 963 691
rect 885 679 889 683
rect 893 679 897 683
rect 901 679 905 683
rect 909 679 913 683
rect 939 679 943 683
rect 947 679 951 683
rect 955 679 959 683
rect 681 639 687 643
rect 683 631 687 635
rect 681 623 687 627
rect 780 626 800 630
rect 806 626 828 630
rect 780 618 798 622
rect 252 536 310 540
rect 360 536 364 540
rect 368 536 372 540
rect 415 536 419 584
rect 423 578 427 582
rect 423 570 427 574
rect 423 562 427 566
rect 423 554 427 558
rect 423 546 427 550
rect 423 538 427 542
rect 254 528 258 532
rect 262 528 266 532
rect 270 528 274 532
rect 278 528 282 532
rect 296 528 300 532
rect 304 528 308 532
rect 360 528 364 532
rect 368 528 372 532
rect 681 560 687 564
rect 683 552 687 556
rect 755 560 761 564
rect 780 563 800 567
rect 806 563 828 567
rect 755 552 759 556
rect 780 555 798 559
rect 813 555 828 559
rect 681 544 687 548
rect 755 544 761 548
rect 780 547 800 551
rect 806 547 828 551
rect 780 539 798 543
rect -21 456 -17 512
rect -13 506 -9 510
rect -13 498 -9 502
rect -13 490 -9 494
rect -13 482 -9 486
rect -13 474 -9 478
rect -13 466 -9 470
rect -13 458 -9 462
rect 156 503 163 507
rect 156 495 160 499
rect 204 498 209 502
rect 156 487 163 491
rect 196 490 209 494
rect 84 480 91 484
rect 415 481 419 505
rect 423 499 427 503
rect 423 491 427 495
rect 423 483 427 487
rect 87 472 91 476
rect 681 513 687 517
rect 683 505 687 509
rect 755 513 761 517
rect 755 505 759 509
rect 813 508 828 512
rect 681 497 687 501
rect 755 497 761 501
rect 780 500 800 504
rect 806 500 828 504
rect 755 489 759 493
rect 780 492 798 496
rect 813 492 828 496
rect 755 481 761 485
rect 806 484 828 488
rect 84 464 91 468
rect 181 467 192 471
rect 181 459 189 463
rect -21 409 -17 425
rect -13 419 -9 423
rect -13 411 -9 415
rect 1 352 5 357
rect 17 352 21 357
rect 25 342 29 357
rect 25 325 29 338
rect 437 397 441 415
rect 453 397 457 415
rect 33 352 37 357
rect 49 352 53 357
rect 33 332 37 337
rect 57 342 61 357
rect 57 325 61 338
rect 286 358 290 368
rect 65 352 69 357
rect 65 332 69 337
rect 31 308 35 312
rect 63 308 67 312
rect 334 358 338 368
rect 461 388 465 415
rect 461 356 465 382
rect 469 397 473 415
rect 485 397 489 415
rect 469 363 473 382
rect 493 388 497 415
rect 493 356 497 382
rect 501 397 505 415
rect 501 363 505 382
rect 509 388 513 415
rect 509 356 513 382
rect 517 397 521 415
rect 517 363 521 382
rect 525 388 529 415
rect 525 356 529 382
rect 533 397 537 415
rect 533 363 537 382
rect 541 388 545 415
rect 541 356 545 382
rect 549 397 553 415
rect 549 363 553 382
rect 557 388 561 415
rect 557 356 561 382
rect 565 397 569 415
rect 565 363 569 382
rect 573 388 577 415
rect 573 356 577 382
rect 581 397 585 415
rect 581 363 585 382
rect 589 388 593 415
rect 589 356 593 382
rect 597 397 601 415
rect 597 363 601 382
rect 605 388 609 415
rect 605 356 609 382
rect 613 397 617 415
rect 613 363 617 382
rect 621 388 625 415
rect 621 356 625 382
rect 629 397 633 415
rect 629 363 633 382
rect 637 388 641 415
rect 637 356 641 382
rect 645 397 649 415
rect 645 363 649 382
rect 653 388 657 415
rect 653 356 657 382
rect 661 397 665 415
rect 939 406 943 428
rect 661 363 665 382
rect 278 338 282 348
rect 302 338 306 348
rect 326 338 330 348
rect 350 338 354 348
rect 468 339 472 343
rect 499 339 503 343
rect 515 339 519 343
rect 531 339 535 343
rect 547 339 551 343
rect 564 339 568 343
rect 580 339 584 343
rect 595 339 599 343
rect 611 339 615 343
rect 627 339 631 343
rect 643 339 647 343
rect 659 339 663 343
rect 1025 406 1029 428
rect 901 375 905 396
rect 955 375 959 396
rect 1011 375 1015 396
rect 1064 397 1068 416
rect 1041 375 1045 396
rect 901 336 905 360
rect 955 336 959 360
rect 1011 336 1015 360
rect 1041 336 1045 360
rect 1072 388 1076 416
rect 1072 356 1076 382
rect 1080 397 1084 416
rect 1080 363 1084 382
rect 1078 339 1082 343
rect 278 312 282 324
rect 326 312 330 324
rect 467 326 473 330
rect 499 326 506 330
rect 515 326 522 330
rect 531 326 538 330
rect 547 326 554 330
rect 563 326 570 330
rect 579 326 586 330
rect 595 326 602 330
rect 611 326 618 330
rect 627 326 634 330
rect 643 326 650 330
rect 659 326 666 330
rect 31 295 38 299
rect 63 295 70 299
rect 262 296 266 308
rect 310 296 314 308
rect 468 307 472 311
rect 499 307 503 311
rect 516 307 520 311
rect 531 307 535 311
rect 547 307 551 311
rect 563 307 567 311
rect 579 307 583 311
rect 595 307 599 311
rect 611 307 615 311
rect 627 307 631 311
rect 643 307 647 311
rect 659 307 663 311
rect 885 310 889 332
rect 467 294 473 298
rect 499 294 506 298
rect 515 294 522 298
rect 531 294 538 298
rect 547 294 554 298
rect 563 294 570 298
rect 579 294 586 298
rect 595 294 602 298
rect 611 294 618 298
rect 627 294 634 298
rect 643 294 650 298
rect 659 294 666 298
rect 955 310 959 332
rect 995 310 999 332
rect 1041 310 1045 332
rect 1078 326 1084 330
rect 1078 308 1082 312
rect 1078 297 1084 301
<< psubstratepdiff >>
rect 228 442 381 443
rect 250 438 367 442
rect 371 438 377 442
<< psubstratepcontact >>
rect 853 708 857 712
rect 439 689 667 693
rect 918 663 922 667
rect 964 663 968 667
rect 853 658 857 662
rect 918 647 922 651
rect 964 647 968 651
rect 918 631 922 635
rect 964 631 968 635
rect 853 626 857 630
rect 3 538 71 542
rect 439 592 443 596
rect 455 592 459 596
rect 471 592 475 596
rect 487 592 491 596
rect 503 592 507 596
rect 519 592 523 596
rect 535 592 539 596
rect 551 592 555 596
rect 567 592 571 596
rect 583 592 587 596
rect 599 592 603 596
rect 615 592 619 596
rect 631 592 635 596
rect 647 592 651 596
rect 858 597 881 601
rect 663 592 667 596
rect 918 584 922 619
rect 964 584 968 619
rect 717 576 721 580
rect 853 579 857 583
rect 918 568 922 572
rect 964 568 968 572
rect 1001 570 1005 574
rect 853 563 857 567
rect 918 552 922 556
rect 964 552 968 556
rect 853 547 857 551
rect 120 503 124 507
rect 227 490 231 494
rect 120 480 124 484
rect 439 513 443 517
rect 455 513 459 517
rect 367 472 371 476
rect 471 513 475 517
rect 487 513 491 517
rect 503 513 507 517
rect 519 513 523 517
rect 535 513 539 517
rect 551 513 555 517
rect 567 513 571 517
rect 583 513 587 517
rect 599 513 603 517
rect 615 513 619 517
rect 631 513 635 517
rect 647 513 651 517
rect 858 518 881 522
rect 663 513 667 517
rect 918 505 922 540
rect 964 505 968 540
rect 1001 538 1005 542
rect 853 500 857 504
rect 918 489 922 493
rect 964 489 968 493
rect 717 481 721 485
rect 853 484 857 488
rect 853 473 861 477
rect 227 467 231 471
rect 885 468 889 472
rect 901 468 905 472
rect 939 468 943 472
rect 367 456 371 460
rect 377 456 381 460
rect 3 433 7 437
rect 19 433 23 437
rect 35 433 39 437
rect 51 433 55 437
rect 228 438 250 442
rect 367 438 371 442
rect 377 438 381 442
rect 67 433 71 437
rect 367 425 371 429
rect 377 425 381 429
rect 367 409 371 413
rect 377 409 381 413
rect 227 401 235 405
rect 262 396 266 400
rect 278 396 282 400
rect 286 396 290 400
rect 302 396 306 400
rect 310 396 314 400
rect 326 396 330 400
rect 334 396 338 400
rect 25 377 29 381
rect 350 396 354 400
rect 461 443 465 447
rect 57 377 61 381
rect 493 443 497 447
rect 509 443 513 447
rect 525 443 529 447
rect 541 443 545 447
rect 557 443 561 447
rect 573 443 577 447
rect 589 443 593 447
rect 605 443 609 447
rect 621 443 625 447
rect 637 443 641 447
rect 955 468 959 472
rect 995 468 999 472
rect 1011 468 1015 472
rect 1025 468 1029 472
rect 1041 468 1045 472
rect 653 443 657 447
rect 1072 443 1076 447
rect 22 281 26 285
rect 38 281 42 285
rect 54 281 58 285
rect 70 281 74 285
rect 442 278 446 282
rect 458 278 462 282
rect 474 278 478 282
rect 490 278 494 282
rect 506 278 510 282
rect 522 278 526 282
rect 538 278 542 282
rect 554 278 558 282
rect 570 278 574 282
rect 586 278 590 282
rect 602 278 606 282
rect 618 278 622 282
rect 634 278 638 282
rect 650 278 654 282
rect 666 278 670 282
rect 262 264 266 268
rect 278 264 282 268
rect 310 264 314 268
rect 326 264 330 268
rect 885 264 889 268
rect 901 264 905 268
rect 1069 281 1073 285
rect 1085 281 1089 285
rect 955 264 959 268
rect 995 264 999 268
rect 1011 264 1015 268
rect 1041 264 1045 268
<< nsubstratencontact >>
rect 762 721 766 725
rect 762 705 766 709
rect 801 708 805 712
rect 883 692 963 696
rect 411 615 415 663
rect 676 655 680 659
rect 762 655 766 659
rect 676 639 680 643
rect 676 623 680 627
rect 801 626 805 630
rect 252 541 310 545
rect 410 536 414 584
rect 676 560 680 564
rect 762 560 766 564
rect 801 563 805 567
rect 676 544 680 548
rect 762 544 766 548
rect 801 547 805 551
rect -26 456 -22 512
rect 163 503 167 507
rect 163 487 167 491
rect 192 490 196 494
rect 80 480 84 484
rect 410 481 414 505
rect 676 513 680 517
rect 762 513 766 517
rect 676 497 680 501
rect 762 497 766 501
rect 801 500 805 504
rect 762 481 766 485
rect 801 484 805 488
rect 80 464 84 468
rect 192 467 196 471
rect -26 409 -22 425
rect 25 338 29 342
rect 57 338 61 342
rect 262 334 266 338
rect 367 358 371 368
rect 461 383 465 387
rect 493 383 497 387
rect 509 383 513 387
rect 525 383 529 387
rect 541 383 545 387
rect 557 383 561 387
rect 573 383 577 387
rect 589 383 593 387
rect 605 383 609 387
rect 621 383 625 387
rect 637 383 641 387
rect 653 383 657 387
rect 918 406 922 428
rect 885 370 889 374
rect 278 334 282 338
rect 286 334 290 338
rect 302 334 306 338
rect 310 334 314 338
rect 326 334 330 338
rect 334 334 338 338
rect 350 334 354 338
rect 901 370 905 374
rect 917 370 921 374
rect 939 370 943 374
rect 955 370 959 374
rect 995 370 999 374
rect 1011 370 1015 374
rect 1025 370 1029 374
rect 1041 370 1045 374
rect 1072 383 1076 387
rect 442 326 446 330
rect 458 326 462 330
rect 474 326 478 330
rect 490 326 494 330
rect 506 326 510 330
rect 522 326 526 330
rect 538 326 542 330
rect 554 326 558 330
rect 570 326 574 330
rect 586 326 590 330
rect 602 326 606 330
rect 618 326 622 330
rect 634 326 638 330
rect 650 326 654 330
rect 666 326 670 330
rect 22 295 26 299
rect 38 295 42 299
rect 54 295 58 299
rect 70 295 74 299
rect 367 296 371 307
rect 442 294 446 298
rect 458 294 462 298
rect 474 294 478 298
rect 490 294 494 298
rect 506 294 510 298
rect 522 294 526 298
rect 538 294 542 298
rect 554 294 558 298
rect 570 294 574 298
rect 586 294 590 298
rect 602 294 606 298
rect 618 294 622 298
rect 634 294 638 298
rect 650 294 654 298
rect 666 294 670 298
rect 918 310 922 331
rect 1069 326 1073 330
rect 1085 326 1089 330
rect 1069 295 1073 299
rect 1085 295 1089 299
<< polysilicon >>
rect 710 718 739 720
rect 743 718 755 720
rect 759 718 761 720
rect 777 713 808 715
rect 828 713 840 715
rect 850 713 852 715
rect 728 710 731 712
rect 735 710 755 712
rect 759 710 761 712
rect 880 710 881 712
rect 878 684 885 686
rect 889 684 893 686
rect 897 684 901 686
rect 905 684 909 686
rect 913 684 939 686
rect 943 684 947 686
rect 951 684 955 686
rect 959 684 966 686
rect 443 675 449 680
rect 443 674 444 675
rect 448 674 449 675
rect 459 675 464 680
rect 459 674 460 675
rect 468 675 472 680
rect 476 675 480 680
rect 484 675 488 680
rect 492 675 496 680
rect 500 675 504 680
rect 508 675 512 680
rect 516 675 520 680
rect 524 675 528 680
rect 532 675 536 680
rect 540 675 544 680
rect 548 675 552 680
rect 556 675 560 680
rect 564 675 568 680
rect 572 675 576 680
rect 580 675 584 680
rect 588 675 592 680
rect 596 675 600 680
rect 604 675 608 680
rect 612 675 616 680
rect 620 675 624 680
rect 628 675 632 680
rect 636 675 640 680
rect 644 675 648 680
rect 652 675 656 680
rect 660 675 664 680
rect 920 683 924 684
rect 420 608 422 666
rect 444 608 446 671
rect 460 608 462 671
rect 468 608 470 671
rect 476 608 478 671
rect 484 608 486 671
rect 492 608 494 671
rect 500 608 502 671
rect 508 608 510 671
rect 516 608 518 671
rect 524 608 526 671
rect 532 608 534 671
rect 540 608 542 671
rect 548 608 550 671
rect 556 608 558 671
rect 564 608 566 671
rect 572 608 574 671
rect 580 608 582 671
rect 588 608 590 671
rect 596 608 598 671
rect 604 608 606 671
rect 612 608 614 671
rect 620 608 622 671
rect 628 608 630 671
rect 636 608 638 671
rect 644 608 646 671
rect 652 608 654 671
rect 660 608 662 671
rect 881 652 885 654
rect 889 652 925 654
rect 929 652 971 654
rect 929 650 934 652
rect 881 644 901 646
rect 905 644 909 646
rect 913 644 925 646
rect 929 644 971 646
rect 929 642 934 644
rect 681 636 683 638
rect 687 636 699 638
rect 703 636 706 638
rect 673 628 683 630
rect 687 628 710 630
rect 714 628 716 630
rect 673 619 675 628
rect 777 623 778 625
rect 798 623 860 625
rect 870 623 872 625
rect 880 620 925 622
rect 417 603 423 608
rect 417 602 418 603
rect 422 602 423 603
rect 443 603 449 608
rect 443 602 444 603
rect 247 533 254 535
rect 258 533 262 535
rect 266 533 270 535
rect 274 533 278 535
rect 282 533 296 535
rect 300 533 304 535
rect 308 533 360 535
rect 364 533 368 535
rect 372 533 379 535
rect 420 582 422 599
rect 448 602 449 603
rect 459 603 464 608
rect 459 602 460 603
rect 468 603 472 608
rect 476 603 480 608
rect 484 603 488 608
rect 492 603 496 608
rect 500 603 504 608
rect 508 603 512 608
rect 516 603 520 608
rect 524 603 528 608
rect 532 603 536 608
rect 540 603 544 608
rect 548 603 552 608
rect 556 603 560 608
rect 564 603 568 608
rect 572 603 576 608
rect 580 603 584 608
rect 588 603 592 608
rect 596 603 600 608
rect 604 603 608 608
rect 612 603 616 608
rect 620 603 624 608
rect 628 603 632 608
rect 636 603 640 608
rect 644 603 648 608
rect 652 603 656 608
rect 660 603 664 608
rect 444 582 446 599
rect 420 574 422 578
rect 444 574 446 578
rect 420 566 422 570
rect 444 566 446 570
rect 420 558 422 562
rect 444 558 446 562
rect 420 550 422 554
rect 444 550 446 554
rect 420 542 422 546
rect 444 542 446 546
rect 284 532 293 533
rect 284 528 289 532
rect 420 529 422 538
rect 444 529 446 538
rect 460 529 462 599
rect 468 529 470 599
rect 476 582 478 599
rect 476 574 478 578
rect 476 529 478 570
rect 484 558 486 599
rect 484 529 486 554
rect 492 550 494 599
rect 500 574 502 599
rect 492 529 494 546
rect 500 529 502 570
rect 508 529 510 599
rect 516 582 518 599
rect 516 529 518 578
rect 524 529 526 599
rect 532 542 534 599
rect 540 582 542 599
rect 540 574 542 578
rect 532 529 534 538
rect 540 529 542 570
rect 548 566 550 599
rect 548 529 550 562
rect 556 529 558 599
rect 564 529 566 599
rect 572 529 574 599
rect 580 529 582 599
rect 588 529 590 599
rect 596 566 598 599
rect 604 574 606 599
rect 612 582 614 599
rect 596 558 598 562
rect 596 550 598 554
rect 596 542 598 546
rect 596 529 598 538
rect 604 529 606 570
rect 612 529 614 578
rect 620 542 622 599
rect 628 566 630 599
rect 628 558 630 562
rect 628 550 630 554
rect 620 529 622 538
rect 628 529 630 546
rect 636 529 638 599
rect 644 566 646 599
rect 652 566 654 599
rect 644 558 646 562
rect 652 558 654 562
rect 644 550 646 554
rect 652 550 654 554
rect 644 542 646 546
rect 644 529 646 538
rect 652 529 654 546
rect 660 542 662 599
rect 929 620 939 622
rect 943 620 947 622
rect 951 620 971 622
rect 929 618 934 620
rect 880 581 925 583
rect 929 581 939 583
rect 943 581 947 583
rect 951 581 971 583
rect 929 579 934 581
rect 880 573 925 575
rect 935 573 939 575
rect 943 573 947 575
rect 951 573 971 575
rect 673 565 716 567
rect 728 565 761 567
rect 673 556 675 565
rect 681 557 683 559
rect 687 557 699 559
rect 703 557 706 559
rect 996 567 1008 569
rect 880 565 885 567
rect 889 565 925 567
rect 777 560 778 562
rect 798 560 860 562
rect 870 560 872 562
rect 929 565 971 567
rect 929 563 934 565
rect 1012 567 1018 569
rect 1012 565 1017 567
rect 710 557 739 559
rect 743 557 755 559
rect 759 557 761 559
rect 673 549 683 551
rect 687 549 710 551
rect 714 549 716 551
rect 880 557 885 559
rect 889 557 925 559
rect 777 552 808 554
rect 828 552 840 554
rect 850 552 852 554
rect 929 557 971 559
rect 929 555 934 557
rect 728 549 731 551
rect 735 549 755 551
rect 759 549 761 551
rect 673 540 675 549
rect 880 549 885 551
rect 889 549 924 551
rect 934 549 971 551
rect 777 544 778 546
rect 798 544 860 546
rect 870 544 872 546
rect 996 543 1008 545
rect 880 541 901 543
rect 905 541 909 543
rect 913 541 925 543
rect 660 529 662 538
rect 284 527 290 528
rect 417 524 423 529
rect 417 523 418 524
rect 422 523 423 524
rect 444 524 448 529
rect -16 510 -14 515
rect -16 502 -14 506
rect -16 494 -14 498
rect -16 486 -14 490
rect -16 478 -14 482
rect -16 470 -14 474
rect -16 462 -14 466
rect -16 449 -14 458
rect 8 449 10 520
rect 16 510 18 512
rect 24 510 26 520
rect 16 502 18 506
rect 24 502 26 506
rect 16 494 18 498
rect 24 494 26 498
rect 16 486 18 490
rect 24 486 26 490
rect 16 478 18 482
rect 24 478 26 482
rect 16 470 18 474
rect 16 462 18 466
rect 16 456 18 458
rect 24 449 26 474
rect 32 470 34 520
rect 40 470 42 520
rect 48 502 50 520
rect 48 494 50 498
rect 48 486 50 490
rect 48 478 50 482
rect 32 456 34 466
rect 40 449 42 466
rect 48 462 50 474
rect 56 470 58 520
rect 64 510 66 520
rect 56 462 58 466
rect 48 449 50 458
rect 56 456 58 458
rect 64 449 66 506
rect 112 500 134 502
rect 138 500 156 502
rect 160 500 162 502
rect 169 498 175 499
rect 169 494 174 498
rect 178 495 199 497
rect 209 495 219 497
rect 224 495 226 497
rect 131 492 142 494
rect 146 492 156 494
rect 160 492 162 494
rect 169 493 175 494
rect 249 492 250 494
rect 85 477 87 479
rect 91 477 108 479
rect 420 503 422 520
rect 460 524 464 529
rect 468 524 472 529
rect 476 524 480 529
rect 484 524 488 529
rect 492 524 496 529
rect 500 524 504 529
rect 508 524 512 529
rect 516 524 520 529
rect 524 524 528 529
rect 532 524 536 529
rect 540 524 544 529
rect 548 524 552 529
rect 556 524 560 529
rect 564 524 568 529
rect 572 524 576 529
rect 580 524 584 529
rect 588 524 592 529
rect 596 524 600 529
rect 604 524 608 529
rect 612 524 616 529
rect 620 524 624 529
rect 628 524 632 529
rect 636 524 640 529
rect 644 524 648 529
rect 652 524 656 529
rect 660 524 664 529
rect 444 503 446 520
rect 420 495 422 499
rect 444 495 446 499
rect 420 487 422 491
rect 444 487 446 491
rect 112 477 113 479
rect 117 477 119 479
rect 420 478 422 483
rect 444 473 446 483
rect 460 473 462 520
rect 468 473 470 520
rect 476 481 478 520
rect 484 473 486 520
rect 492 473 494 520
rect 500 473 502 520
rect 508 473 510 520
rect 516 473 518 520
rect 524 473 526 520
rect 532 473 534 520
rect 540 473 542 520
rect 548 473 550 520
rect 556 473 558 520
rect 564 473 566 520
rect 572 473 574 520
rect 580 473 582 520
rect 588 495 590 520
rect 588 473 590 491
rect 596 487 598 520
rect 596 473 598 483
rect 604 473 606 520
rect 612 473 614 520
rect 620 473 622 520
rect 628 503 630 520
rect 636 503 638 520
rect 628 495 630 499
rect 628 487 630 491
rect 628 473 630 483
rect 636 473 638 499
rect 644 487 646 520
rect 644 473 646 483
rect 652 473 654 520
rect 660 503 662 520
rect 681 510 683 512
rect 687 510 699 512
rect 703 510 706 512
rect 710 510 739 512
rect 743 510 755 512
rect 759 510 761 512
rect 673 502 683 504
rect 687 502 710 504
rect 714 502 716 504
rect 777 505 808 507
rect 828 505 840 507
rect 850 505 852 507
rect 929 541 971 543
rect 929 539 934 541
rect 1012 543 1018 545
rect 728 502 731 504
rect 735 502 755 504
rect 759 502 761 504
rect 660 495 662 499
rect 673 493 675 502
rect 880 502 885 504
rect 889 502 925 504
rect 777 497 778 499
rect 798 497 860 499
rect 870 497 872 499
rect 929 502 971 504
rect 929 500 934 502
rect 710 494 739 496
rect 743 494 755 496
rect 759 494 761 496
rect 660 487 662 491
rect 880 494 885 496
rect 889 494 925 496
rect 777 489 808 491
rect 828 489 840 491
rect 850 489 852 491
rect 929 494 971 496
rect 929 492 934 494
rect 728 486 731 488
rect 735 486 755 488
rect 759 486 761 488
rect 660 473 662 483
rect 880 486 893 488
rect 897 486 925 488
rect 929 486 955 488
rect 959 486 971 488
rect 929 484 934 486
rect 951 475 954 477
rect 1037 475 1040 477
rect 77 469 87 471
rect 91 469 101 471
rect 105 469 107 471
rect 77 460 79 469
rect 169 467 175 468
rect 250 469 262 471
rect 362 469 372 471
rect 169 463 174 467
rect 178 464 179 466
rect 189 464 234 466
rect 239 464 241 466
rect 169 462 175 463
rect 249 461 262 463
rect 362 461 372 463
rect -16 423 -14 440
rect 8 423 10 440
rect 16 423 18 444
rect -16 415 -14 419
rect 8 415 10 419
rect -16 406 -14 411
rect 8 401 10 411
rect 16 409 18 419
rect 24 401 26 440
rect 32 401 34 444
rect 40 409 42 440
rect 48 409 50 440
rect 56 401 58 444
rect 64 423 66 440
rect 250 422 254 424
rect 258 422 310 424
rect 314 422 350 424
rect 354 422 358 424
rect 362 422 384 424
rect 64 415 66 419
rect 250 414 254 416
rect 258 414 270 416
rect 274 414 278 416
rect 282 414 286 416
rect 290 414 294 416
rect 298 414 302 416
rect 306 414 310 416
rect 314 414 318 416
rect 322 414 326 416
rect 330 414 334 416
rect 338 414 342 416
rect 346 414 358 416
rect 362 414 384 416
rect 64 401 66 411
rect 298 403 301 405
rect 346 403 349 405
rect 30 391 32 393
rect 62 391 64 393
rect 299 393 301 403
rect 22 374 24 376
rect 22 357 24 367
rect 22 322 24 345
rect 30 335 32 384
rect 347 393 349 403
rect 450 390 452 465
rect 466 463 468 465
rect 498 463 500 465
rect 514 463 516 465
rect 530 463 532 465
rect 546 463 548 465
rect 562 463 564 465
rect 578 463 580 465
rect 594 463 596 465
rect 610 463 612 465
rect 626 463 628 465
rect 642 463 644 465
rect 658 463 660 465
rect 458 440 460 442
rect 458 415 460 427
rect 291 384 293 385
rect 54 374 56 376
rect 54 357 56 367
rect 30 322 32 323
rect 54 322 56 345
rect 62 335 64 384
rect 291 376 293 378
rect 291 368 293 370
rect 291 355 293 356
rect 62 322 64 323
rect 22 320 23 322
rect 30 319 31 322
rect 54 320 55 322
rect 62 319 63 322
rect 267 308 269 351
rect 299 353 301 387
rect 347 353 349 387
rect 458 353 460 390
rect 466 380 468 450
rect 490 440 492 442
rect 490 415 492 427
rect 466 353 468 354
rect 490 353 492 390
rect 498 380 500 450
rect 506 440 508 442
rect 506 415 508 427
rect 498 353 500 354
rect 506 353 508 390
rect 514 380 516 450
rect 522 440 524 442
rect 522 415 524 427
rect 514 353 516 354
rect 522 353 524 390
rect 530 380 532 450
rect 538 440 540 442
rect 538 415 540 427
rect 530 353 532 354
rect 538 353 540 390
rect 546 380 548 450
rect 554 440 556 442
rect 554 415 556 427
rect 546 353 548 354
rect 554 353 556 390
rect 562 380 564 450
rect 570 440 572 442
rect 570 415 572 427
rect 562 353 564 354
rect 570 353 572 390
rect 578 380 580 450
rect 586 440 588 442
rect 586 415 588 427
rect 578 353 580 354
rect 586 353 588 390
rect 594 380 596 450
rect 602 440 604 442
rect 602 415 604 427
rect 594 353 596 354
rect 602 353 604 390
rect 610 380 612 450
rect 618 440 620 442
rect 618 415 620 427
rect 610 353 612 354
rect 618 353 620 390
rect 626 380 628 450
rect 634 440 636 442
rect 634 415 636 427
rect 626 353 628 354
rect 634 353 636 390
rect 642 380 644 450
rect 952 465 954 475
rect 1038 465 1040 475
rect 1071 473 1073 481
rect 1079 473 1081 481
rect 1077 463 1079 465
rect 944 450 946 451
rect 650 440 652 442
rect 650 415 652 427
rect 642 353 644 354
rect 650 353 652 390
rect 658 380 660 450
rect 944 436 946 440
rect 944 428 946 430
rect 944 403 946 404
rect 658 353 660 354
rect 299 339 301 341
rect 347 339 349 341
rect 465 337 467 338
rect 462 336 467 337
rect 471 336 473 338
rect 496 337 499 338
rect 493 336 499 337
rect 503 336 505 338
rect 512 336 515 338
rect 519 336 521 338
rect 528 336 531 338
rect 535 336 537 338
rect 544 336 547 338
rect 551 336 553 338
rect 561 337 563 338
rect 558 336 563 337
rect 567 336 569 338
rect 577 337 579 338
rect 574 336 579 337
rect 583 336 585 338
rect 592 336 595 338
rect 599 336 601 338
rect 608 336 611 338
rect 615 336 617 338
rect 624 336 627 338
rect 631 336 633 338
rect 640 336 643 338
rect 647 336 649 338
rect 656 336 659 338
rect 663 336 665 338
rect 464 331 467 333
rect 471 331 473 333
rect 496 331 499 333
rect 503 331 505 333
rect 512 331 515 333
rect 519 331 521 333
rect 528 331 531 333
rect 535 331 537 333
rect 544 331 547 333
rect 551 331 553 333
rect 560 331 563 333
rect 567 331 569 333
rect 576 331 579 333
rect 583 331 585 333
rect 592 331 595 333
rect 599 331 601 333
rect 608 331 611 333
rect 615 331 617 333
rect 624 331 627 333
rect 631 331 633 333
rect 640 331 643 333
rect 647 331 649 333
rect 656 331 659 333
rect 663 331 665 333
rect 890 332 892 399
rect 952 401 954 453
rect 1038 401 1040 453
rect 1069 440 1071 442
rect 1069 416 1071 428
rect 952 375 954 377
rect 1038 375 1040 377
rect 898 360 900 363
rect 1008 360 1010 363
rect 1069 353 1071 390
rect 1077 380 1079 450
rect 1077 353 1079 354
rect 275 324 277 327
rect 323 324 325 327
rect 464 323 466 331
rect 496 323 498 331
rect 512 323 514 331
rect 528 323 530 331
rect 544 323 546 331
rect 560 323 562 331
rect 576 323 578 331
rect 592 323 594 331
rect 608 323 610 331
rect 624 323 626 331
rect 640 323 642 331
rect 656 323 658 331
rect 60 305 63 307
rect 67 305 69 307
rect 28 300 31 302
rect 35 300 37 302
rect 60 300 63 302
rect 67 300 69 302
rect 28 293 30 300
rect 60 293 62 300
rect 267 294 269 296
rect 28 292 37 293
rect 32 288 37 292
rect 28 287 37 288
rect 60 292 69 293
rect 64 288 69 292
rect 60 287 69 288
rect 28 280 30 287
rect 60 280 62 287
rect 267 286 269 288
rect 28 278 31 280
rect 35 278 37 280
rect 60 278 63 280
rect 67 278 69 280
rect 267 279 269 280
rect 275 277 277 312
rect 323 277 325 312
rect 465 305 467 306
rect 462 304 467 305
rect 471 304 473 306
rect 496 304 499 306
rect 503 304 505 306
rect 513 305 515 306
rect 510 304 515 305
rect 519 304 521 306
rect 528 304 531 306
rect 535 304 537 306
rect 544 304 547 306
rect 551 304 553 306
rect 560 304 563 306
rect 567 304 569 306
rect 576 304 579 306
rect 583 304 585 306
rect 592 304 595 306
rect 599 304 601 306
rect 608 304 611 306
rect 615 304 617 306
rect 624 304 627 306
rect 631 304 633 306
rect 640 304 643 306
rect 647 304 649 306
rect 890 306 892 310
rect 656 304 659 306
rect 663 304 665 306
rect 464 299 467 301
rect 471 299 473 301
rect 496 299 499 301
rect 503 299 505 301
rect 512 299 515 301
rect 519 299 521 301
rect 528 299 531 301
rect 535 299 537 301
rect 544 299 547 301
rect 551 299 553 301
rect 560 299 563 301
rect 567 299 569 301
rect 576 299 579 301
rect 583 299 585 301
rect 592 299 595 301
rect 599 299 601 301
rect 608 299 611 301
rect 615 299 617 301
rect 624 299 627 301
rect 631 299 633 301
rect 640 299 643 301
rect 647 299 649 301
rect 656 299 659 301
rect 663 299 665 301
rect 464 289 466 299
rect 496 289 498 299
rect 512 289 514 299
rect 528 289 530 299
rect 544 289 546 299
rect 560 289 562 299
rect 576 289 578 299
rect 592 289 594 299
rect 608 289 610 299
rect 624 289 626 299
rect 640 289 642 299
rect 656 289 658 299
rect 890 298 892 300
rect 890 285 892 286
rect 464 277 466 285
rect 496 277 498 285
rect 512 277 514 285
rect 528 277 530 285
rect 544 277 546 285
rect 560 277 562 285
rect 576 277 578 285
rect 592 277 594 285
rect 608 277 610 285
rect 624 277 626 285
rect 640 277 642 285
rect 656 277 658 285
rect 898 283 900 336
rect 1008 283 1010 336
rect 1075 331 1078 333
rect 1082 331 1084 333
rect 1075 323 1077 331
rect 1075 302 1078 304
rect 1082 302 1084 304
rect 1075 292 1077 302
rect 60 271 63 272
rect 58 270 63 271
rect 67 270 69 272
rect 275 269 277 271
rect 464 275 467 277
rect 471 275 473 277
rect 496 275 499 277
rect 503 275 505 277
rect 512 275 515 277
rect 519 275 521 277
rect 528 275 531 277
rect 535 275 537 277
rect 544 275 547 277
rect 551 275 553 277
rect 560 275 563 277
rect 567 275 569 277
rect 576 275 579 277
rect 583 275 585 277
rect 592 275 595 277
rect 599 275 601 277
rect 608 275 611 277
rect 615 275 617 277
rect 624 275 627 277
rect 631 275 633 277
rect 640 275 643 277
rect 647 275 649 277
rect 656 275 659 277
rect 663 275 665 277
rect 323 269 325 271
rect 463 271 467 272
rect 465 270 467 271
rect 471 270 473 272
rect 496 270 499 272
rect 503 270 505 272
rect 511 271 515 272
rect 513 270 515 271
rect 519 270 521 272
rect 528 270 531 272
rect 535 270 537 272
rect 544 270 547 272
rect 551 270 553 272
rect 560 270 563 272
rect 567 270 569 272
rect 576 270 579 272
rect 583 270 585 272
rect 592 270 595 272
rect 599 270 601 272
rect 608 270 611 272
rect 615 270 617 272
rect 624 270 627 272
rect 631 270 633 272
rect 640 270 643 272
rect 647 270 649 272
rect 656 270 659 272
rect 663 270 665 272
rect 898 269 900 271
rect 1075 280 1077 288
rect 1075 278 1078 280
rect 1082 278 1084 280
rect 1008 269 1010 271
<< polycontact >>
rect 706 717 710 721
rect 724 710 728 714
rect 773 712 777 716
rect 876 708 880 712
rect 966 684 970 688
rect 876 680 880 684
rect 444 671 448 675
rect 460 671 464 675
rect 468 671 472 675
rect 476 671 480 675
rect 484 671 488 675
rect 492 671 496 675
rect 500 671 504 675
rect 508 671 512 675
rect 516 671 520 675
rect 524 671 528 675
rect 532 671 536 675
rect 540 671 544 675
rect 548 671 552 675
rect 556 671 560 675
rect 564 671 568 675
rect 572 671 576 675
rect 580 671 584 675
rect 588 671 592 675
rect 596 671 600 675
rect 604 671 608 675
rect 612 671 616 675
rect 620 671 624 675
rect 628 671 632 675
rect 636 671 640 675
rect 644 671 648 675
rect 652 671 656 675
rect 920 679 924 683
rect 660 671 664 675
rect 418 666 422 670
rect 925 650 929 654
rect 971 650 975 654
rect 925 642 929 646
rect 971 642 975 646
rect 706 635 710 639
rect 669 618 673 622
rect 773 622 777 626
rect 876 618 880 622
rect 418 599 422 603
rect 379 533 383 537
rect 444 599 448 603
rect 460 599 464 603
rect 468 599 472 603
rect 476 599 480 603
rect 484 599 488 603
rect 492 599 496 603
rect 500 599 504 603
rect 508 599 512 603
rect 516 599 520 603
rect 524 599 528 603
rect 532 599 536 603
rect 540 599 544 603
rect 548 599 552 603
rect 556 599 560 603
rect 564 599 568 603
rect 572 599 576 603
rect 580 599 584 603
rect 588 599 592 603
rect 596 599 600 603
rect 604 599 608 603
rect 612 599 616 603
rect 620 599 624 603
rect 628 599 632 603
rect 636 599 640 603
rect 644 599 648 603
rect 652 599 656 603
rect 660 599 664 603
rect 245 529 249 533
rect 289 528 293 532
rect 925 618 929 622
rect 971 618 975 622
rect 925 579 929 583
rect 971 579 975 583
rect 724 565 728 569
rect 971 571 975 575
rect 669 555 673 559
rect 706 556 710 560
rect 876 563 880 567
rect 773 559 777 563
rect 925 563 929 567
rect 971 563 975 567
rect 1008 565 1012 569
rect 724 549 728 553
rect 773 551 777 555
rect 876 555 880 559
rect 925 555 929 559
rect 971 555 975 559
rect 669 538 673 542
rect 876 547 880 551
rect 773 543 777 547
rect 971 547 975 551
rect 876 539 880 543
rect 8 520 12 524
rect 24 520 28 524
rect 32 520 36 524
rect 40 520 44 524
rect 48 520 52 524
rect 56 520 60 524
rect 64 520 68 524
rect 418 520 422 524
rect -18 515 -14 519
rect 108 500 112 504
rect 127 492 131 496
rect 174 494 178 498
rect 245 490 249 494
rect 108 477 112 481
rect 444 520 448 524
rect 460 520 464 524
rect 468 520 472 524
rect 476 520 480 524
rect 484 520 488 524
rect 492 520 496 524
rect 500 520 504 524
rect 508 520 512 524
rect 516 520 520 524
rect 524 520 528 524
rect 532 520 536 524
rect 540 520 544 524
rect 548 520 552 524
rect 556 520 560 524
rect 564 520 568 524
rect 572 520 576 524
rect 580 520 584 524
rect 588 520 592 524
rect 596 520 600 524
rect 604 520 608 524
rect 612 520 616 524
rect 620 520 624 524
rect 628 520 632 524
rect 636 520 640 524
rect 644 520 648 524
rect 652 520 656 524
rect 660 520 664 524
rect 418 474 422 478
rect 706 509 710 513
rect 724 502 728 506
rect 773 504 777 508
rect 925 539 929 543
rect 971 539 975 543
rect 1008 541 1012 545
rect 669 491 673 495
rect 706 493 710 497
rect 876 500 880 504
rect 773 496 777 500
rect 925 500 929 504
rect 971 500 975 504
rect 724 486 728 490
rect 773 488 777 492
rect 876 492 880 496
rect 925 492 929 496
rect 971 492 975 496
rect 876 484 880 488
rect 925 484 929 488
rect 971 484 975 488
rect 947 475 951 479
rect 1033 475 1037 479
rect 73 458 77 462
rect 444 469 448 473
rect 460 469 464 473
rect 468 469 472 473
rect 484 469 488 473
rect 492 469 496 473
rect 500 469 504 473
rect 508 469 512 473
rect 516 469 520 473
rect 524 469 528 473
rect 532 469 536 473
rect 540 469 544 473
rect 548 469 552 473
rect 556 469 560 473
rect 564 469 568 473
rect 572 469 576 473
rect 580 469 584 473
rect 588 469 592 473
rect 596 469 600 473
rect 604 469 608 473
rect 612 469 616 473
rect 620 469 624 473
rect 628 469 632 473
rect 636 469 640 473
rect 644 469 648 473
rect 652 469 656 473
rect 660 469 664 473
rect 174 463 178 467
rect 245 459 249 463
rect -18 440 -14 444
rect 8 440 12 444
rect 24 440 28 444
rect -18 402 -14 406
rect 40 440 44 444
rect 48 440 52 444
rect 64 440 68 444
rect 384 420 388 424
rect 384 412 388 416
rect 294 403 298 407
rect 342 403 346 407
rect 8 397 12 401
rect 24 397 28 401
rect 32 397 36 401
rect 56 397 60 401
rect 64 397 68 401
rect 290 385 294 389
rect 266 351 270 355
rect 23 318 27 322
rect 31 318 35 322
rect 55 318 59 322
rect 63 318 67 322
rect 56 305 60 309
rect 290 351 294 355
rect 943 451 947 455
rect 1071 469 1075 473
rect 1079 469 1083 473
rect 889 399 893 403
rect 458 349 462 353
rect 466 349 470 353
rect 490 349 494 353
rect 498 349 502 353
rect 506 349 510 353
rect 514 349 518 353
rect 522 349 526 353
rect 530 349 534 353
rect 538 349 542 353
rect 546 349 550 353
rect 554 349 558 353
rect 562 349 566 353
rect 570 349 574 353
rect 578 349 582 353
rect 586 349 590 353
rect 594 349 598 353
rect 602 349 606 353
rect 610 349 614 353
rect 618 349 622 353
rect 626 349 630 353
rect 634 349 638 353
rect 642 349 646 353
rect 650 349 654 353
rect 658 349 662 353
rect 461 337 465 341
rect 492 337 496 341
rect 508 336 512 340
rect 524 336 528 340
rect 540 336 544 340
rect 557 337 561 341
rect 573 337 577 341
rect 588 336 592 340
rect 604 336 608 340
rect 620 336 624 340
rect 636 336 640 340
rect 652 336 656 340
rect 943 399 947 403
rect 898 363 902 367
rect 1008 363 1012 367
rect 1069 349 1073 353
rect 1077 349 1081 353
rect 275 327 279 331
rect 323 327 327 331
rect 463 319 467 323
rect 495 319 499 323
rect 511 319 515 323
rect 527 319 531 323
rect 543 319 547 323
rect 559 319 563 323
rect 575 319 579 323
rect 591 319 595 323
rect 607 319 611 323
rect 623 319 627 323
rect 639 319 643 323
rect 655 319 659 323
rect 28 288 32 292
rect 60 288 64 292
rect 56 271 60 275
rect 266 275 270 279
rect 461 305 465 309
rect 492 304 496 308
rect 509 305 513 309
rect 524 304 528 308
rect 540 304 544 308
rect 556 304 560 308
rect 572 304 576 308
rect 588 304 592 308
rect 604 304 608 308
rect 620 304 624 308
rect 636 304 640 308
rect 652 304 656 308
rect 463 285 467 289
rect 495 285 499 289
rect 511 285 515 289
rect 527 285 531 289
rect 543 285 547 289
rect 559 285 563 289
rect 575 285 579 289
rect 591 285 595 289
rect 607 285 611 289
rect 623 285 627 289
rect 639 285 643 289
rect 655 285 659 289
rect 889 281 893 285
rect 1074 319 1078 323
rect 1074 288 1078 292
rect 461 267 465 271
rect 492 268 496 272
rect 509 267 513 271
rect 524 268 528 272
rect 540 268 544 272
rect 556 268 560 272
rect 572 268 576 272
rect 588 268 592 272
rect 604 268 608 272
rect 620 268 624 272
rect 636 268 640 272
rect 652 268 656 272
<< metal1 >>
rect 667 707 668 711
rect 676 705 680 725
rect 707 721 710 725
rect 707 705 710 717
rect 717 705 721 725
rect 724 709 728 710
rect 731 709 735 725
rect 743 721 749 724
rect 761 721 762 725
rect 746 717 749 721
rect 750 714 755 717
rect 762 709 766 721
rect 806 712 810 725
rect 828 717 840 720
rect 831 712 834 717
rect 853 712 857 725
rect 761 705 762 709
rect 805 708 806 712
rect 852 708 853 712
rect 875 708 876 712
rect 806 705 810 708
rect 853 705 857 708
rect 426 689 439 693
rect 667 689 857 695
rect 883 691 963 692
rect 426 687 667 689
rect 426 679 430 687
rect 418 670 422 671
rect 440 665 447 668
rect 451 665 463 668
rect 467 665 479 668
rect 483 665 495 668
rect 499 665 511 668
rect 515 665 527 668
rect 531 665 543 668
rect 547 665 559 668
rect 563 665 575 668
rect 579 665 591 668
rect 595 665 607 668
rect 611 665 623 668
rect 627 665 639 668
rect 643 665 655 668
rect 659 665 663 668
rect 427 657 439 660
rect 443 657 455 660
rect 459 657 503 660
rect 507 657 551 660
rect 555 657 599 660
rect 603 657 615 660
rect 619 657 647 660
rect 651 657 663 660
rect 667 657 668 661
rect 676 659 680 669
rect 707 655 710 667
rect 717 655 721 689
rect 724 659 728 660
rect 731 659 735 689
rect 762 678 846 682
rect 746 667 749 669
rect 750 664 755 667
rect 762 659 766 678
rect 806 665 810 678
rect 853 673 857 689
rect 880 687 883 691
rect 872 680 876 683
rect 966 683 970 684
rect 853 669 876 673
rect 853 662 857 669
rect 743 655 749 658
rect 853 655 857 658
rect 885 651 888 679
rect 680 639 681 643
rect 691 639 699 642
rect 707 639 710 643
rect 676 627 680 639
rect 691 635 694 639
rect 687 632 690 635
rect 680 623 681 627
rect 667 620 669 621
rect 427 617 439 620
rect 443 617 471 620
rect 475 617 535 620
rect 539 617 567 620
rect 571 617 615 620
rect 619 618 669 620
rect 619 617 670 618
rect 411 584 415 615
rect 440 611 447 614
rect 451 611 463 614
rect 467 611 479 614
rect 483 611 495 614
rect 499 611 511 614
rect 515 611 527 614
rect 531 611 543 614
rect 547 611 559 614
rect 563 611 575 614
rect 579 611 591 614
rect 595 611 607 614
rect 611 611 623 614
rect 627 611 639 614
rect 643 611 655 614
rect 659 611 663 614
rect 430 592 439 596
rect 443 592 455 596
rect 459 592 471 596
rect 475 592 487 596
rect 491 592 503 596
rect 507 592 519 596
rect 523 592 535 596
rect 539 592 551 596
rect 555 592 567 596
rect 571 592 583 596
rect 587 592 599 596
rect 603 592 615 596
rect 619 592 631 596
rect 635 592 647 596
rect 651 592 663 596
rect 440 586 447 589
rect 451 586 463 589
rect 467 586 479 589
rect 483 586 495 589
rect 499 586 511 589
rect 515 586 527 589
rect 531 586 543 589
rect 547 586 559 589
rect 563 586 575 589
rect 579 586 591 589
rect 595 586 607 589
rect 611 586 623 589
rect 627 586 639 589
rect 643 586 655 589
rect 659 586 663 589
rect -10 538 3 542
rect 71 538 231 544
rect 252 540 310 541
rect -10 536 71 538
rect -10 528 -6 536
rect -18 519 -14 520
rect 4 514 11 517
rect 15 514 27 517
rect 31 514 35 517
rect 39 514 43 517
rect 47 514 59 517
rect 63 514 67 517
rect -22 456 -21 512
rect -9 506 19 509
rect 23 506 67 509
rect 120 507 124 538
rect -9 498 19 501
rect 23 498 51 501
rect 55 498 71 501
rect -9 490 19 493
rect 23 490 51 493
rect 55 490 67 493
rect 71 489 72 493
rect -9 482 19 485
rect 23 482 51 485
rect 55 482 71 485
rect 80 484 84 507
rect 109 504 112 507
rect 109 481 112 500
rect 120 484 124 503
rect 134 507 138 538
rect 163 527 220 531
rect 163 507 167 527
rect 127 491 131 492
rect -9 474 19 477
rect 23 474 51 477
rect 55 474 71 477
rect -9 466 19 469
rect 23 466 35 469
rect 39 466 51 469
rect 55 466 71 469
rect 80 468 84 480
rect 91 472 94 475
rect 95 468 98 472
rect 95 465 101 468
rect -9 458 19 461
rect 23 458 51 461
rect 55 458 67 461
rect 71 458 73 462
rect -25 425 -21 456
rect 4 452 11 455
rect 19 452 27 455
rect 35 452 43 455
rect 47 452 51 455
rect 63 452 67 455
rect -6 433 3 437
rect 7 433 19 437
rect 23 433 35 437
rect 39 433 51 437
rect 55 433 67 437
rect 4 427 11 430
rect 15 427 27 430
rect 31 427 43 430
rect 47 427 51 430
rect 55 427 59 430
rect 63 427 67 430
rect -22 409 -21 425
rect -9 419 3 422
rect 7 419 19 422
rect 23 419 67 422
rect -9 411 3 414
rect 7 411 67 414
rect 80 409 84 464
rect -25 329 -21 409
rect 4 404 11 407
rect 15 404 27 407
rect 31 404 43 407
rect 47 404 59 407
rect 63 405 76 407
rect 80 405 90 409
rect 109 405 112 477
rect 63 404 73 405
rect -18 401 -14 402
rect -25 299 -21 325
rect -17 307 -14 397
rect 8 396 12 397
rect 25 396 29 397
rect 33 396 37 397
rect 57 396 61 397
rect 65 396 69 397
rect 33 391 37 392
rect 65 391 69 392
rect 75 381 79 393
rect -6 377 25 381
rect 29 377 57 381
rect 61 377 79 381
rect 82 389 90 405
rect 82 385 86 389
rect -10 285 -6 377
rect 1 363 4 367
rect 17 363 20 367
rect 1 360 6 363
rect 17 360 25 363
rect 33 363 36 367
rect 49 363 52 367
rect 33 360 37 363
rect 49 360 57 363
rect 65 363 68 367
rect 65 360 69 363
rect 1 357 4 360
rect 17 357 20 360
rect 33 357 36 360
rect 49 357 52 360
rect 65 357 68 360
rect 12 345 25 349
rect 29 345 57 349
rect 82 349 90 385
rect 61 345 90 349
rect 3 325 25 329
rect 33 337 37 338
rect 29 325 57 329
rect 65 337 69 338
rect 82 329 90 345
rect 61 325 90 329
rect 82 324 90 325
rect 23 317 27 318
rect 31 317 35 318
rect 55 317 59 318
rect 63 317 67 318
rect 31 312 35 313
rect 63 312 67 313
rect 82 320 86 324
rect 3 303 75 305
rect 0 302 75 303
rect 82 299 90 320
rect 3 295 22 299
rect 26 295 31 299
rect 42 295 54 299
rect 58 295 63 299
rect 74 295 90 299
rect -10 281 22 285
rect 26 281 31 285
rect 42 281 54 285
rect 58 281 63 285
rect 28 273 31 276
rect 41 275 75 278
rect 60 265 63 268
rect 82 264 90 295
rect 94 278 97 401
rect 120 397 124 480
rect 134 397 138 503
rect 153 495 156 498
rect 149 491 152 495
rect 163 491 167 503
rect 197 494 201 527
rect 227 522 231 538
rect 249 536 252 540
rect 310 536 360 540
rect 364 536 368 540
rect 414 536 415 584
rect 427 578 439 581
rect 443 578 471 581
rect 475 578 519 581
rect 523 578 535 581
rect 539 578 615 581
rect 667 581 672 582
rect 619 578 672 581
rect 676 580 680 623
rect 707 576 710 635
rect 717 580 721 643
rect 724 576 728 581
rect 731 580 735 643
rect 762 580 766 643
rect 806 630 810 643
rect 853 630 857 643
rect 800 626 801 630
rect 805 626 806 630
rect 852 626 853 630
rect 857 626 858 630
rect 798 618 799 622
rect 806 583 810 626
rect 853 601 857 626
rect 870 618 871 622
rect 875 618 876 622
rect 857 597 858 601
rect 853 583 857 597
rect 871 579 876 583
rect 427 570 439 573
rect 443 570 471 573
rect 475 570 503 573
rect 507 570 535 573
rect 539 570 599 573
rect 603 570 667 573
rect 427 562 439 565
rect 443 562 551 565
rect 555 562 599 565
rect 603 562 631 565
rect 635 562 647 565
rect 667 565 668 566
rect 651 562 668 565
rect 676 564 680 576
rect 680 560 681 564
rect 691 560 699 563
rect 707 560 710 572
rect 427 554 439 557
rect 443 554 487 557
rect 491 554 599 557
rect 603 554 631 557
rect 635 554 647 557
rect 667 557 669 558
rect 651 555 669 557
rect 651 554 670 555
rect 427 546 439 549
rect 443 546 487 549
rect 491 546 599 549
rect 603 546 631 549
rect 635 546 647 549
rect 667 549 668 550
rect 651 546 668 549
rect 676 548 680 560
rect 691 556 694 560
rect 687 553 690 556
rect 680 544 681 548
rect 427 538 439 541
rect 443 538 535 541
rect 539 538 599 541
rect 603 538 615 541
rect 619 538 647 541
rect 651 538 663 541
rect 667 538 669 542
rect 241 529 245 532
rect 379 532 383 533
rect 227 518 245 522
rect 209 499 219 502
rect 212 494 215 499
rect 227 494 231 518
rect 146 488 152 491
rect 244 490 245 494
rect 163 389 167 487
rect 197 471 201 490
rect 196 467 201 471
rect 189 459 190 463
rect 197 389 201 467
rect 227 471 231 490
rect 227 442 231 467
rect 239 459 240 463
rect 244 459 245 463
rect 227 438 228 442
rect 227 409 231 438
rect 254 429 257 528
rect 254 413 257 425
rect 262 409 265 528
rect 270 413 273 528
rect 278 413 281 528
rect 287 516 291 518
rect 296 516 299 528
rect 304 516 307 528
rect 360 516 363 528
rect 368 516 371 528
rect 286 413 289 476
rect 294 413 297 476
rect 302 413 305 476
rect 310 429 313 476
rect 310 413 313 425
rect 318 413 321 476
rect 326 413 329 476
rect 334 413 337 476
rect 342 413 345 476
rect 350 429 353 476
rect 358 429 361 476
rect 367 468 371 472
rect 367 460 371 464
rect 367 442 371 456
rect 367 429 371 438
rect 350 409 353 425
rect 358 413 361 425
rect 367 421 371 425
rect 367 413 371 417
rect 377 460 381 518
rect 411 505 415 536
rect 440 532 447 535
rect 451 532 463 535
rect 467 532 479 535
rect 483 532 495 535
rect 499 532 511 535
rect 515 532 527 535
rect 531 532 543 535
rect 547 532 559 535
rect 563 532 575 535
rect 579 532 591 535
rect 595 532 607 535
rect 611 532 623 535
rect 627 532 639 535
rect 643 532 655 535
rect 659 532 663 535
rect 676 517 680 544
rect 430 513 439 517
rect 443 513 455 517
rect 459 513 471 517
rect 475 513 487 517
rect 491 513 503 517
rect 507 513 519 517
rect 523 513 535 517
rect 539 513 551 517
rect 555 513 567 517
rect 571 513 583 517
rect 587 513 599 517
rect 603 513 615 517
rect 619 513 631 517
rect 635 513 647 517
rect 651 513 663 517
rect 680 513 681 517
rect 691 513 699 516
rect 707 513 710 556
rect 440 507 447 510
rect 451 507 463 510
rect 467 507 479 510
rect 483 507 495 510
rect 499 507 511 510
rect 515 507 527 510
rect 531 507 543 510
rect 547 507 559 510
rect 563 507 575 510
rect 579 507 591 510
rect 595 507 607 510
rect 611 507 623 510
rect 627 507 639 510
rect 643 507 655 510
rect 659 507 663 510
rect 414 481 415 505
rect 427 499 439 502
rect 443 499 631 502
rect 635 499 663 502
rect 667 499 668 503
rect 676 501 680 513
rect 691 509 694 513
rect 687 506 690 509
rect 680 497 681 501
rect 707 497 710 509
rect 427 491 439 494
rect 443 491 583 494
rect 587 491 631 494
rect 635 491 663 494
rect 667 491 669 495
rect 427 483 439 486
rect 443 483 599 486
rect 603 483 631 486
rect 635 483 647 486
rect 651 483 663 486
rect 667 483 668 487
rect 676 481 680 497
rect 377 442 381 456
rect 377 429 381 438
rect 377 421 381 425
rect 388 420 389 424
rect 377 413 381 417
rect 388 412 389 416
rect 227 405 235 409
rect 262 407 266 409
rect 294 407 298 409
rect 310 407 314 409
rect 342 407 346 409
rect 220 389 223 401
rect 227 400 235 401
rect 227 397 262 400
rect 231 396 262 397
rect 266 396 278 400
rect 282 396 286 400
rect 290 396 302 400
rect 306 396 310 400
rect 314 396 326 400
rect 330 396 334 400
rect 338 396 350 400
rect 354 396 372 400
rect 231 393 235 396
rect 94 264 97 274
rect 102 264 105 302
rect 212 264 215 351
rect 220 278 223 385
rect 220 264 223 274
rect 227 268 235 393
rect 250 385 290 388
rect 294 385 306 388
rect 350 385 372 388
rect 286 375 289 378
rect 334 375 337 378
rect 286 368 289 371
rect 334 368 337 371
rect 367 368 371 369
rect 411 360 415 481
rect 440 476 447 479
rect 451 476 463 479
rect 467 476 479 479
rect 483 476 495 479
rect 499 476 511 479
rect 515 476 527 479
rect 531 476 543 479
rect 547 476 559 479
rect 563 476 575 479
rect 579 476 591 479
rect 595 476 607 479
rect 611 476 623 479
rect 627 476 639 479
rect 643 476 655 479
rect 659 476 673 479
rect 676 477 685 481
rect 418 473 422 474
rect 670 469 673 476
rect 250 351 266 354
rect 270 351 290 354
rect 294 351 306 354
rect 350 351 372 354
rect 246 334 262 338
rect 266 334 278 338
rect 282 334 286 338
rect 290 334 302 338
rect 306 334 310 338
rect 314 334 326 338
rect 330 334 334 338
rect 338 334 350 338
rect 354 334 372 338
rect 246 324 250 334
rect 274 327 275 331
rect 322 327 323 331
rect 411 330 415 356
rect 419 338 422 469
rect 445 468 449 469
rect 461 468 465 469
rect 469 468 473 469
rect 469 463 473 464
rect 485 468 489 469
rect 493 468 497 469
rect 501 468 505 469
rect 509 468 513 469
rect 517 468 521 469
rect 525 468 529 469
rect 533 468 537 469
rect 541 468 545 469
rect 549 468 553 469
rect 557 468 561 469
rect 565 468 569 469
rect 573 468 577 469
rect 581 468 585 469
rect 589 468 593 469
rect 597 468 601 469
rect 605 468 609 469
rect 613 468 617 469
rect 621 468 625 469
rect 629 468 633 469
rect 637 468 641 469
rect 645 468 649 469
rect 653 468 657 469
rect 661 468 665 469
rect 485 463 489 464
rect 501 463 505 464
rect 461 447 465 448
rect 517 463 521 464
rect 493 447 497 448
rect 533 463 537 464
rect 509 447 513 448
rect 549 463 553 464
rect 525 447 529 448
rect 565 463 569 464
rect 541 447 545 448
rect 581 463 585 464
rect 557 447 561 448
rect 597 463 601 464
rect 573 447 577 448
rect 613 463 617 464
rect 589 447 593 448
rect 629 463 633 464
rect 605 447 609 448
rect 645 463 649 464
rect 621 447 625 448
rect 661 463 665 464
rect 637 447 641 448
rect 677 461 685 477
rect 707 477 710 493
rect 717 485 721 576
rect 724 564 728 565
rect 731 564 735 576
rect 762 564 766 576
rect 798 571 803 575
rect 806 567 810 579
rect 828 572 840 575
rect 831 567 834 572
rect 853 567 857 579
rect 870 571 876 575
rect 885 572 888 647
rect 893 635 896 679
rect 901 667 904 679
rect 909 667 912 679
rect 918 667 922 669
rect 901 651 904 663
rect 909 651 912 663
rect 918 659 922 663
rect 918 651 922 655
rect 743 560 749 563
rect 761 560 762 564
rect 800 563 801 567
rect 805 563 806 567
rect 852 563 853 567
rect 857 563 858 567
rect 875 563 876 567
rect 724 548 728 549
rect 731 548 735 560
rect 746 556 749 560
rect 750 553 755 556
rect 762 548 766 560
rect 798 555 799 559
rect 806 551 810 563
rect 828 556 840 559
rect 831 551 834 556
rect 853 551 857 563
rect 870 555 871 559
rect 875 555 876 559
rect 885 556 888 568
rect 761 544 762 548
rect 800 547 801 551
rect 805 547 806 551
rect 852 547 853 551
rect 857 547 858 551
rect 875 547 876 551
rect 724 501 728 502
rect 731 501 735 544
rect 762 517 766 544
rect 798 539 799 543
rect 743 513 749 516
rect 761 513 762 517
rect 746 509 749 513
rect 750 506 755 509
rect 762 501 766 513
rect 806 504 810 547
rect 853 522 857 547
rect 870 539 871 543
rect 875 539 876 543
rect 857 518 858 522
rect 828 509 840 512
rect 831 504 834 509
rect 853 504 857 518
rect 885 509 888 552
rect 743 497 749 500
rect 761 497 762 501
rect 800 500 801 504
rect 805 500 806 504
rect 852 500 853 504
rect 857 500 858 504
rect 875 500 876 504
rect 724 485 728 486
rect 731 485 735 497
rect 746 493 749 497
rect 750 490 755 493
rect 762 485 766 497
rect 798 492 799 496
rect 806 488 810 500
rect 828 493 840 496
rect 831 488 834 493
rect 853 488 857 500
rect 870 492 871 496
rect 875 492 876 496
rect 885 493 888 505
rect 893 493 896 631
rect 901 540 904 647
rect 909 540 912 647
rect 918 643 922 647
rect 918 635 922 639
rect 918 627 922 631
rect 918 619 922 623
rect 939 619 942 679
rect 947 619 950 679
rect 955 635 958 679
rect 964 667 968 669
rect 964 659 968 663
rect 964 651 968 655
rect 975 650 976 654
rect 964 643 968 647
rect 975 642 976 646
rect 964 635 968 639
rect 922 597 923 601
rect 918 580 922 584
rect 939 588 942 615
rect 947 588 950 615
rect 918 572 922 576
rect 918 564 922 568
rect 939 572 942 584
rect 947 572 950 584
rect 918 556 922 560
rect 918 548 922 552
rect 918 540 922 544
rect 761 481 762 485
rect 805 484 806 488
rect 852 484 853 488
rect 875 484 876 488
rect 717 469 721 481
rect 677 457 681 461
rect 653 447 657 448
rect 250 320 278 324
rect 282 320 326 324
rect 330 320 372 324
rect 367 307 371 320
rect 419 306 422 334
rect 430 443 461 447
rect 465 443 477 447
rect 485 443 493 447
rect 497 443 509 447
rect 513 443 525 447
rect 529 443 541 447
rect 545 443 557 447
rect 561 443 573 447
rect 577 443 589 447
rect 593 443 605 447
rect 609 443 621 447
rect 625 443 637 447
rect 641 443 653 447
rect 657 443 670 447
rect 262 293 265 296
rect 310 293 313 296
rect 367 293 371 296
rect 262 286 265 289
rect 310 286 313 289
rect 426 282 430 443
rect 461 442 465 443
rect 493 442 497 443
rect 509 442 513 443
rect 525 442 529 443
rect 541 442 545 443
rect 557 442 561 443
rect 573 442 577 443
rect 589 442 593 443
rect 605 442 609 443
rect 621 442 625 443
rect 637 442 641 443
rect 653 442 657 443
rect 437 422 440 427
rect 437 419 445 422
rect 453 422 456 427
rect 453 419 461 422
rect 437 415 440 419
rect 453 415 456 419
rect 469 415 472 427
rect 485 422 488 427
rect 485 419 493 422
rect 501 422 504 427
rect 501 419 509 422
rect 517 422 520 427
rect 517 419 525 422
rect 533 422 536 427
rect 533 419 541 422
rect 549 422 552 427
rect 549 419 557 422
rect 565 422 568 427
rect 565 419 573 422
rect 581 422 584 427
rect 581 419 589 422
rect 597 422 600 427
rect 597 419 605 422
rect 613 422 616 427
rect 613 419 621 422
rect 629 422 632 427
rect 629 419 637 422
rect 645 422 648 427
rect 645 419 653 422
rect 661 422 664 427
rect 661 419 665 422
rect 485 415 488 419
rect 501 415 504 419
rect 517 415 520 419
rect 533 415 536 419
rect 549 415 552 419
rect 565 415 568 419
rect 581 415 584 419
rect 597 415 600 419
rect 613 415 616 419
rect 629 415 632 419
rect 645 415 648 419
rect 661 415 664 419
rect 439 390 445 394
rect 449 390 461 394
rect 465 390 477 394
rect 485 390 493 394
rect 461 387 465 388
rect 497 390 509 394
rect 493 387 497 388
rect 513 390 525 394
rect 509 387 513 388
rect 529 390 541 394
rect 525 387 529 388
rect 545 390 557 394
rect 541 387 545 388
rect 561 390 573 394
rect 557 387 561 388
rect 577 390 589 394
rect 573 387 577 388
rect 593 390 605 394
rect 589 387 593 388
rect 609 390 621 394
rect 605 387 609 388
rect 625 390 637 394
rect 621 387 625 388
rect 641 390 653 394
rect 637 387 641 388
rect 677 394 685 457
rect 657 390 685 394
rect 653 387 657 388
rect 461 382 465 383
rect 439 356 445 360
rect 449 356 461 360
rect 469 382 473 383
rect 493 382 497 383
rect 465 356 477 360
rect 490 356 493 360
rect 501 382 505 383
rect 509 382 513 383
rect 497 356 509 360
rect 517 382 521 383
rect 525 382 529 383
rect 513 356 525 360
rect 533 382 537 383
rect 541 382 545 383
rect 529 356 541 360
rect 549 382 553 383
rect 557 382 561 383
rect 545 356 557 360
rect 565 382 569 383
rect 573 382 577 383
rect 561 356 573 360
rect 581 382 585 383
rect 589 382 593 383
rect 577 356 589 360
rect 597 382 601 383
rect 605 382 609 383
rect 593 356 605 360
rect 613 382 617 383
rect 621 382 625 383
rect 609 356 621 360
rect 629 382 633 383
rect 637 382 641 383
rect 625 356 637 360
rect 645 382 649 383
rect 653 382 657 383
rect 641 356 653 360
rect 661 382 665 383
rect 677 360 685 390
rect 657 356 681 360
rect 451 348 455 349
rect 459 348 463 349
rect 467 348 471 349
rect 491 348 495 349
rect 499 348 503 349
rect 507 348 511 349
rect 515 348 519 349
rect 523 348 527 349
rect 531 348 535 349
rect 539 348 543 349
rect 547 348 551 349
rect 555 348 559 349
rect 563 348 567 349
rect 571 348 575 349
rect 579 348 583 349
rect 587 348 591 349
rect 595 348 599 349
rect 603 348 607 349
rect 611 348 615 349
rect 619 348 623 349
rect 627 348 631 349
rect 635 348 639 349
rect 643 348 647 349
rect 651 348 655 349
rect 659 348 663 349
rect 451 343 455 344
rect 468 343 471 344
rect 499 343 503 344
rect 461 336 465 337
rect 515 343 519 344
rect 492 336 496 337
rect 531 343 535 344
rect 547 343 551 344
rect 564 343 567 344
rect 580 343 583 344
rect 595 343 599 344
rect 557 336 561 337
rect 573 336 577 337
rect 611 343 615 344
rect 627 343 631 344
rect 643 343 647 344
rect 659 343 663 344
rect 439 334 477 336
rect 436 333 477 334
rect 490 333 670 336
rect 677 330 685 356
rect 439 326 442 330
rect 446 326 451 330
rect 455 326 458 330
rect 462 326 467 330
rect 473 326 474 330
rect 494 326 499 330
rect 510 326 515 330
rect 526 326 531 330
rect 542 326 547 330
rect 558 326 563 330
rect 574 326 579 330
rect 590 326 595 330
rect 606 326 611 330
rect 622 326 627 330
rect 638 326 643 330
rect 654 326 659 330
rect 670 326 685 330
rect 467 319 468 323
rect 499 319 500 323
rect 515 319 516 323
rect 531 319 532 323
rect 547 319 548 323
rect 563 319 564 323
rect 579 319 580 323
rect 595 319 596 323
rect 611 319 612 323
rect 627 319 628 323
rect 643 319 644 323
rect 659 319 660 323
rect 448 312 455 315
rect 464 312 471 315
rect 496 312 503 315
rect 512 312 519 315
rect 528 312 535 315
rect 544 312 551 315
rect 560 312 567 315
rect 576 312 583 315
rect 592 312 599 315
rect 608 312 615 315
rect 624 312 631 315
rect 640 312 647 315
rect 656 312 663 315
rect 468 311 471 312
rect 499 311 503 312
rect 461 304 465 305
rect 516 311 519 312
rect 531 311 535 312
rect 509 304 513 305
rect 547 311 551 312
rect 563 311 567 312
rect 579 311 583 312
rect 595 311 599 312
rect 611 311 615 312
rect 627 311 631 312
rect 643 311 647 312
rect 659 311 663 312
rect 439 302 477 304
rect 436 301 477 302
rect 490 301 670 304
rect 677 298 685 326
rect 439 294 442 298
rect 446 294 451 298
rect 455 294 458 298
rect 462 294 467 298
rect 473 294 474 298
rect 494 294 499 298
rect 510 294 515 298
rect 526 294 531 298
rect 542 294 547 298
rect 558 294 563 298
rect 574 294 579 298
rect 590 294 595 298
rect 606 294 611 298
rect 622 294 627 298
rect 638 294 643 298
rect 654 294 659 298
rect 670 294 685 298
rect 467 285 468 289
rect 499 285 500 289
rect 515 285 516 289
rect 531 285 532 289
rect 547 285 548 289
rect 563 285 564 289
rect 579 285 580 289
rect 595 285 596 289
rect 611 285 612 289
rect 627 285 628 289
rect 643 285 644 289
rect 659 285 660 289
rect 250 275 266 278
rect 426 278 442 282
rect 446 278 451 282
rect 455 278 458 282
rect 462 278 467 282
rect 473 278 474 282
rect 494 278 499 282
rect 510 278 515 282
rect 526 278 531 282
rect 542 278 547 282
rect 558 278 563 282
rect 574 278 579 282
rect 590 278 595 282
rect 606 278 611 282
rect 622 278 627 282
rect 638 278 643 282
rect 654 278 659 282
rect 270 275 306 278
rect 350 275 372 278
rect 439 272 477 275
rect 490 272 670 275
rect 461 271 465 272
rect 227 264 262 268
rect 266 264 278 268
rect 282 264 310 268
rect 314 264 326 268
rect 330 264 372 268
rect 509 271 513 272
rect 468 264 471 265
rect 448 261 454 264
rect 464 261 471 264
rect 496 262 502 265
rect 516 264 519 265
rect 512 261 519 264
rect 528 262 534 265
rect 544 262 550 265
rect 560 262 566 265
rect 576 262 582 265
rect 592 262 598 265
rect 608 262 614 265
rect 624 262 630 265
rect 640 262 646 265
rect 656 262 662 265
rect 677 261 685 294
rect 731 469 735 481
rect 689 275 692 465
rect 717 447 721 465
rect 762 461 766 481
rect 806 461 810 484
rect 853 481 857 484
rect 885 481 888 489
rect 893 481 896 489
rect 901 481 904 536
rect 909 481 912 536
rect 922 518 923 522
rect 918 501 922 505
rect 918 493 922 497
rect 918 485 922 489
rect 939 481 942 568
rect 947 481 950 568
rect 955 493 958 631
rect 964 627 968 631
rect 964 619 968 623
rect 975 618 976 622
rect 968 597 969 601
rect 964 580 968 584
rect 975 579 976 583
rect 964 572 968 576
rect 975 571 976 575
rect 964 564 968 568
rect 975 563 976 567
rect 1001 566 1005 570
rect 964 556 968 560
rect 975 555 976 559
rect 964 548 968 552
rect 975 547 976 551
rect 964 540 968 544
rect 975 539 976 543
rect 1001 542 1005 546
rect 968 518 969 522
rect 964 501 968 505
rect 975 500 976 504
rect 964 493 968 497
rect 975 492 976 496
rect 955 481 958 489
rect 964 485 968 489
rect 975 484 976 488
rect 853 477 861 481
rect 885 479 889 481
rect 947 479 951 481
rect 955 479 959 481
rect 995 479 999 481
rect 1033 479 1037 481
rect 1041 479 1045 481
rect 1064 476 1074 479
rect 1078 476 1089 479
rect 846 455 849 473
rect 853 472 861 473
rect 853 469 885 472
rect 857 468 885 469
rect 889 468 901 472
rect 913 468 939 472
rect 943 468 955 472
rect 991 468 995 472
rect 999 468 1011 472
rect 1029 468 1041 472
rect 857 465 861 468
rect 697 305 700 333
rect 689 261 692 271
rect 697 261 700 301
rect 838 264 841 399
rect 846 284 849 451
rect 846 264 849 280
rect 853 268 861 465
rect 901 467 905 468
rect 955 467 959 468
rect 1011 467 1015 468
rect 1041 467 1045 468
rect 1072 468 1076 469
rect 1080 468 1084 469
rect 1080 463 1084 464
rect 881 451 905 454
rect 913 451 943 454
rect 947 451 959 454
rect 1072 447 1076 448
rect 1064 443 1072 447
rect 1076 443 1088 447
rect 1072 442 1076 443
rect 939 435 942 440
rect 1025 435 1028 440
rect 918 428 922 429
rect 939 428 942 431
rect 1025 428 1028 431
rect 1064 422 1067 428
rect 1064 419 1072 422
rect 1064 416 1067 419
rect 1080 416 1083 428
rect 881 399 889 402
rect 893 399 905 402
rect 913 399 943 402
rect 947 399 959 402
rect 901 374 905 375
rect 955 374 959 375
rect 1011 374 1015 375
rect 1064 390 1072 394
rect 1041 374 1045 375
rect 877 370 885 374
rect 889 370 901 374
rect 913 370 917 374
rect 921 370 939 374
rect 943 370 955 374
rect 991 370 995 374
rect 999 370 1011 374
rect 1029 370 1041 374
rect 1076 390 1088 394
rect 1072 387 1076 388
rect 1072 382 1076 383
rect 877 360 881 370
rect 897 363 898 367
rect 1007 363 1008 367
rect 881 356 901 360
rect 913 356 955 360
rect 918 331 922 356
rect 991 356 1011 360
rect 1025 356 1041 360
rect 1064 356 1072 360
rect 1080 382 1084 383
rect 1076 356 1088 360
rect 1070 348 1074 349
rect 1078 348 1082 349
rect 1078 343 1082 344
rect 885 305 888 310
rect 918 305 922 310
rect 1066 326 1069 330
rect 1073 326 1078 330
rect 1084 326 1085 330
rect 1078 319 1079 323
rect 1075 312 1082 315
rect 955 305 958 310
rect 995 305 998 310
rect 1041 305 1044 310
rect 885 298 888 301
rect 955 298 958 301
rect 995 298 998 301
rect 1041 298 1044 301
rect 1066 295 1069 299
rect 1073 297 1078 299
rect 1084 297 1085 299
rect 1073 295 1085 297
rect 1078 288 1079 292
rect 881 281 889 284
rect 893 281 905 284
rect 913 281 959 284
rect 1066 281 1069 285
rect 1073 281 1078 285
rect 1084 281 1085 285
rect 901 268 905 269
rect 955 268 959 269
rect 1011 268 1015 269
rect 1041 268 1045 269
rect 853 264 885 268
rect 889 264 901 268
rect 913 264 955 268
rect 991 264 995 268
rect 999 264 1011 268
rect 1025 264 1041 268
rect 1075 265 1081 268
<< m2contact >>
rect 668 707 672 711
rect 724 705 728 709
rect 746 713 750 717
rect 769 712 773 716
rect 831 708 835 712
rect 871 708 875 712
rect 426 675 430 679
rect 444 675 448 679
rect 418 671 422 675
rect 460 675 464 679
rect 468 675 472 679
rect 476 675 480 679
rect 484 675 488 679
rect 492 675 496 679
rect 500 675 504 679
rect 508 675 512 679
rect 516 675 520 679
rect 524 675 528 679
rect 532 675 536 679
rect 540 675 544 679
rect 548 675 552 679
rect 556 675 560 679
rect 564 675 568 679
rect 572 675 576 679
rect 580 675 584 679
rect 588 675 592 679
rect 596 675 600 679
rect 604 675 608 679
rect 612 675 616 679
rect 620 675 624 679
rect 628 675 632 679
rect 636 675 640 679
rect 644 675 648 679
rect 652 675 656 679
rect 660 675 664 679
rect 436 664 440 668
rect 668 657 672 661
rect 846 678 850 682
rect 746 663 750 667
rect 769 662 773 666
rect 876 687 880 691
rect 868 679 872 683
rect 916 679 920 683
rect 966 679 970 683
rect 876 669 880 673
rect 724 655 728 659
rect 690 631 694 635
rect 436 610 440 614
rect 418 603 422 607
rect 444 603 448 607
rect 460 603 464 607
rect 468 603 472 607
rect 476 603 480 607
rect 484 603 488 607
rect 492 603 496 607
rect 500 603 504 607
rect 508 603 512 607
rect 516 603 520 607
rect 524 603 528 607
rect 532 603 536 607
rect 540 603 544 607
rect 548 603 552 607
rect 556 603 560 607
rect 564 603 568 607
rect 572 603 576 607
rect 580 603 584 607
rect 588 603 592 607
rect 596 603 600 607
rect 604 603 608 607
rect 612 603 616 607
rect 620 603 624 607
rect 628 603 632 607
rect 636 603 640 607
rect 644 603 648 607
rect 652 603 656 607
rect 660 603 664 607
rect 426 592 430 596
rect 436 585 440 589
rect -10 524 -6 528
rect 8 524 12 528
rect -18 520 -14 524
rect 24 524 28 528
rect 32 524 36 528
rect 40 524 44 528
rect 48 524 52 528
rect 56 524 60 528
rect 64 524 68 528
rect 0 513 4 517
rect 72 489 76 493
rect 220 527 224 531
rect 127 487 131 491
rect 94 472 98 476
rect 0 451 4 455
rect -18 444 -14 448
rect 8 444 12 448
rect 24 444 28 448
rect 40 444 44 448
rect 48 444 52 448
rect 64 444 68 448
rect -10 433 -6 437
rect 0 426 4 430
rect 0 404 4 408
rect 73 401 77 405
rect -18 397 -14 401
rect -25 325 -21 329
rect 8 392 12 396
rect 25 392 29 396
rect 33 392 37 396
rect 57 392 61 396
rect 65 392 69 396
rect 75 393 79 397
rect -18 303 -14 307
rect -10 377 -6 381
rect 86 385 90 389
rect -25 295 -21 299
rect 25 360 29 364
rect 57 360 61 364
rect -1 325 3 329
rect 33 338 37 342
rect 65 338 69 342
rect 23 313 27 317
rect 31 313 35 317
rect 55 313 59 317
rect 63 313 67 317
rect -1 303 3 307
rect 86 320 90 324
rect 75 302 79 306
rect -1 295 3 299
rect 32 288 36 292
rect 64 288 68 292
rect 24 272 28 276
rect 75 274 79 278
rect 56 264 60 268
rect 94 401 98 405
rect 109 401 113 405
rect 120 393 124 397
rect 149 495 153 499
rect 170 494 174 498
rect 245 536 249 540
rect 769 622 773 626
rect 799 618 803 622
rect 871 618 875 622
rect 853 597 857 601
rect 668 562 672 566
rect 668 546 672 550
rect 690 552 694 556
rect 237 528 241 532
rect 285 528 289 532
rect 379 528 383 532
rect 245 518 249 522
rect 212 490 216 494
rect 240 490 244 494
rect 134 393 138 397
rect 170 463 174 467
rect 190 459 194 463
rect 163 385 167 389
rect 240 459 244 463
rect 287 518 291 522
rect 377 518 381 522
rect 436 531 440 535
rect 418 524 422 528
rect 444 524 448 528
rect 460 524 464 528
rect 468 524 472 528
rect 476 524 480 528
rect 484 524 488 528
rect 492 524 496 528
rect 500 524 504 528
rect 508 524 512 528
rect 516 524 520 528
rect 524 524 528 528
rect 532 524 536 528
rect 540 524 544 528
rect 548 524 552 528
rect 556 524 560 528
rect 564 524 568 528
rect 572 524 576 528
rect 580 524 584 528
rect 588 524 592 528
rect 596 524 600 528
rect 604 524 608 528
rect 612 524 616 528
rect 620 524 624 528
rect 628 524 632 528
rect 636 524 640 528
rect 644 524 648 528
rect 652 524 656 528
rect 660 524 664 528
rect 426 513 430 517
rect 436 506 440 510
rect 668 499 672 503
rect 690 505 694 509
rect 668 483 672 487
rect 389 420 393 424
rect 389 412 393 416
rect 197 385 201 389
rect 220 401 224 405
rect 262 403 266 407
rect 310 403 314 407
rect 227 393 231 397
rect 220 385 224 389
rect 212 351 216 355
rect 101 302 105 306
rect 94 274 98 278
rect 220 274 224 278
rect 246 385 250 389
rect 286 371 290 375
rect 334 371 338 375
rect 367 369 371 373
rect 436 476 440 480
rect 418 469 422 473
rect 411 356 415 360
rect 246 351 250 355
rect 270 327 274 331
rect 318 327 322 331
rect 445 464 449 468
rect 461 464 465 468
rect 469 464 473 468
rect 485 464 489 468
rect 493 464 497 468
rect 501 464 505 468
rect 509 464 513 468
rect 517 464 521 468
rect 525 464 529 468
rect 533 464 537 468
rect 541 464 545 468
rect 549 464 553 468
rect 557 464 561 468
rect 565 464 569 468
rect 573 464 577 468
rect 581 464 585 468
rect 589 464 593 468
rect 597 464 601 468
rect 605 464 609 468
rect 613 464 617 468
rect 621 464 625 468
rect 629 464 633 468
rect 637 464 641 468
rect 645 464 649 468
rect 653 464 657 468
rect 661 464 665 468
rect 670 465 674 469
rect 724 560 728 564
rect 918 669 922 673
rect 929 650 933 654
rect 831 563 835 567
rect 871 563 875 567
rect 724 544 728 548
rect 746 552 750 556
rect 769 559 773 563
rect 799 555 803 559
rect 769 551 773 555
rect 871 555 875 559
rect 831 547 835 551
rect 871 547 875 551
rect 724 497 728 501
rect 769 543 773 547
rect 799 539 803 543
rect 746 505 750 509
rect 769 504 773 508
rect 871 539 875 543
rect 853 518 857 522
rect 831 500 835 504
rect 871 500 875 504
rect 724 481 728 485
rect 746 489 750 493
rect 769 496 773 500
rect 799 492 803 496
rect 769 488 773 492
rect 871 492 875 496
rect 929 642 933 646
rect 929 618 933 622
rect 964 669 968 673
rect 976 650 980 654
rect 976 642 980 646
rect 923 597 927 601
rect 929 579 933 583
rect 929 563 933 567
rect 929 555 933 559
rect 831 484 835 488
rect 871 484 875 488
rect 707 473 711 477
rect 681 457 685 461
rect 418 334 422 338
rect 411 326 415 330
rect 246 320 250 324
rect 418 302 422 306
rect 426 443 430 447
rect 670 443 674 447
rect 262 289 266 293
rect 310 289 314 293
rect 367 289 371 293
rect 445 419 449 423
rect 461 419 465 423
rect 493 419 497 423
rect 509 419 513 423
rect 525 419 529 423
rect 541 419 545 423
rect 557 419 561 423
rect 573 419 577 423
rect 589 419 593 423
rect 605 419 609 423
rect 621 419 625 423
rect 637 419 641 423
rect 653 419 657 423
rect 435 356 439 360
rect 469 383 473 387
rect 501 383 505 387
rect 517 383 521 387
rect 533 383 537 387
rect 549 383 553 387
rect 565 383 569 387
rect 581 383 585 387
rect 597 383 601 387
rect 613 383 617 387
rect 629 383 633 387
rect 645 383 649 387
rect 661 383 665 387
rect 681 356 685 360
rect 451 344 455 348
rect 459 344 463 348
rect 467 344 471 348
rect 491 344 495 348
rect 499 344 503 348
rect 507 344 511 348
rect 515 344 519 348
rect 523 344 527 348
rect 531 344 535 348
rect 539 344 543 348
rect 547 344 551 348
rect 555 344 559 348
rect 563 344 567 348
rect 571 344 575 348
rect 579 344 583 348
rect 587 344 591 348
rect 595 344 599 348
rect 603 344 607 348
rect 611 344 615 348
rect 619 344 623 348
rect 627 344 631 348
rect 635 344 639 348
rect 643 344 647 348
rect 651 344 655 348
rect 659 344 663 348
rect 435 334 439 338
rect 670 333 674 337
rect 435 326 439 330
rect 468 319 472 323
rect 500 319 504 323
rect 516 319 520 323
rect 532 319 536 323
rect 548 319 552 323
rect 564 319 568 323
rect 580 319 584 323
rect 596 319 600 323
rect 612 319 616 323
rect 628 319 632 323
rect 644 319 648 323
rect 660 319 664 323
rect 444 312 448 316
rect 460 312 464 316
rect 492 312 496 316
rect 508 312 512 316
rect 524 312 528 316
rect 540 312 544 316
rect 556 312 560 316
rect 572 312 576 316
rect 588 312 592 316
rect 604 312 608 316
rect 620 312 624 316
rect 636 312 640 316
rect 652 312 656 316
rect 435 302 439 306
rect 670 301 674 305
rect 468 285 472 289
rect 500 285 504 289
rect 516 285 520 289
rect 532 285 536 289
rect 548 285 552 289
rect 564 285 568 289
rect 580 285 584 289
rect 596 285 600 289
rect 612 285 616 289
rect 628 285 632 289
rect 644 285 648 289
rect 660 285 664 289
rect 246 274 250 278
rect 670 271 674 275
rect 444 260 448 264
rect 460 260 464 264
rect 492 261 496 265
rect 508 260 512 264
rect 524 261 528 265
rect 540 261 544 265
rect 556 261 560 265
rect 572 261 576 265
rect 588 261 592 265
rect 604 261 608 265
rect 620 261 624 265
rect 636 261 640 265
rect 652 261 656 265
rect 689 465 693 469
rect 717 465 721 469
rect 731 465 735 469
rect 762 457 766 461
rect 929 539 933 543
rect 923 518 927 522
rect 929 500 933 504
rect 929 492 933 496
rect 929 484 933 488
rect 976 618 980 622
rect 969 597 973 601
rect 976 579 980 583
rect 976 571 980 575
rect 976 563 980 567
rect 1012 565 1016 569
rect 976 555 980 559
rect 976 547 980 551
rect 976 539 980 543
rect 1012 541 1016 545
rect 969 518 973 522
rect 976 500 980 504
rect 976 492 980 496
rect 976 484 980 488
rect 806 457 810 461
rect 846 473 850 477
rect 885 475 889 479
rect 955 475 959 479
rect 995 475 999 479
rect 1041 475 1045 479
rect 717 443 721 447
rect 853 465 857 469
rect 846 451 850 455
rect 838 399 842 403
rect 696 333 700 337
rect 696 301 700 305
rect 689 271 693 275
rect 846 280 850 284
rect 1072 464 1076 468
rect 1080 464 1084 468
rect 877 451 881 455
rect 918 429 922 433
rect 939 431 943 435
rect 1025 431 1029 435
rect 1072 419 1076 423
rect 877 399 881 403
rect 893 363 897 367
rect 1003 363 1007 367
rect 877 356 881 360
rect 1080 383 1084 387
rect 1070 344 1074 348
rect 1078 344 1082 348
rect 885 301 889 305
rect 918 301 922 305
rect 1079 319 1083 323
rect 1071 312 1075 316
rect 955 301 959 305
rect 995 301 999 305
rect 1041 301 1045 305
rect 1079 288 1083 292
rect 877 280 881 284
rect 1071 264 1075 268
<< metal2 >>
rect 750 713 769 716
rect 672 709 686 710
rect 672 707 724 709
rect 683 706 724 707
rect 835 709 871 712
rect 875 709 881 712
rect 667 686 834 688
rect 419 685 834 686
rect 419 683 671 685
rect 419 675 422 683
rect 419 607 422 671
rect 71 535 215 537
rect -17 534 215 535
rect -17 532 74 534
rect -17 524 -14 532
rect -17 448 -14 520
rect -17 401 -14 444
rect -10 437 -6 524
rect -10 381 -6 433
rect 0 455 3 513
rect 0 430 3 451
rect 8 448 11 524
rect 16 456 19 512
rect 24 448 27 524
rect 32 456 35 524
rect 40 448 43 524
rect 48 448 51 524
rect 56 456 59 524
rect 64 448 67 524
rect 212 521 215 534
rect 220 536 245 540
rect 220 531 224 536
rect 241 529 285 532
rect 289 529 379 532
rect 419 528 422 603
rect 237 521 240 528
rect 212 518 240 521
rect 249 518 287 522
rect 291 518 377 522
rect 153 495 170 498
rect 76 491 90 492
rect 76 489 127 491
rect 87 488 127 489
rect 216 491 240 494
rect 244 490 250 493
rect 98 472 138 475
rect 419 473 422 524
rect 135 467 138 472
rect 250 468 262 471
rect 362 468 372 471
rect 426 596 430 675
rect 426 517 430 592
rect 135 464 170 467
rect 194 459 240 462
rect 244 460 262 463
rect 362 460 372 463
rect 426 447 430 513
rect 436 614 439 664
rect 436 589 439 610
rect 444 607 447 675
rect 460 607 463 675
rect 468 607 471 675
rect 476 607 479 675
rect 484 607 487 675
rect 492 607 495 675
rect 500 607 503 675
rect 508 607 511 675
rect 516 607 519 675
rect 524 607 527 675
rect 532 607 535 675
rect 540 607 543 675
rect 548 607 551 675
rect 556 607 559 675
rect 564 607 567 675
rect 572 607 575 675
rect 580 607 583 675
rect 588 607 591 675
rect 596 607 599 675
rect 604 607 607 675
rect 612 607 615 675
rect 620 607 623 675
rect 628 607 631 675
rect 636 607 639 675
rect 644 607 647 675
rect 652 607 655 675
rect 660 607 663 675
rect 831 672 834 685
rect 846 687 876 691
rect 846 682 850 687
rect 872 680 916 683
rect 920 680 966 683
rect 868 672 871 679
rect 831 669 871 672
rect 880 669 918 673
rect 922 669 964 673
rect 750 663 769 666
rect 672 659 686 660
rect 672 657 724 659
rect 683 656 724 657
rect 881 651 929 654
rect 933 651 976 654
rect 881 643 929 646
rect 933 643 976 646
rect 694 631 735 634
rect 732 626 735 631
rect 732 623 769 626
rect 803 618 871 621
rect 875 619 929 622
rect 933 619 976 622
rect 436 535 439 585
rect 436 510 439 531
rect 444 528 447 603
rect 460 528 463 603
rect 468 528 471 603
rect 476 528 479 603
rect 484 528 487 603
rect 492 528 495 603
rect 500 528 503 603
rect 508 528 511 603
rect 516 528 519 603
rect 524 528 527 603
rect 532 528 535 603
rect 540 528 543 603
rect 548 528 551 603
rect 556 528 559 603
rect 564 528 567 603
rect 572 528 575 603
rect 580 528 583 603
rect 588 528 591 603
rect 596 528 599 603
rect 604 528 607 603
rect 612 528 615 603
rect 620 528 623 603
rect 628 528 631 603
rect 636 528 639 603
rect 644 528 647 603
rect 652 528 655 603
rect 660 528 663 603
rect 857 597 923 601
rect 927 597 969 601
rect 880 580 929 583
rect 933 580 976 583
rect 880 572 925 575
rect 935 572 976 575
rect 672 564 686 565
rect 672 562 724 564
rect 683 561 724 562
rect 835 564 871 567
rect 875 564 929 567
rect 933 564 976 567
rect 996 566 1012 569
rect 1016 566 1018 569
rect 694 552 735 555
rect 803 555 871 558
rect 875 556 929 559
rect 933 556 976 559
rect 750 552 769 555
rect 672 548 686 549
rect 672 546 724 548
rect 683 545 724 546
rect 732 547 735 552
rect 835 548 871 551
rect 875 548 924 551
rect 934 548 976 551
rect 732 544 769 547
rect 803 539 871 542
rect 875 540 929 543
rect 933 540 976 543
rect 996 542 1012 545
rect 1016 542 1018 545
rect 436 480 439 506
rect 444 475 447 524
rect 460 475 463 524
rect 468 475 471 524
rect 476 481 479 524
rect 484 475 487 524
rect 492 475 495 524
rect 500 475 503 524
rect 508 475 511 524
rect 516 475 519 524
rect 524 475 527 524
rect 532 475 535 524
rect 540 475 543 524
rect 548 475 551 524
rect 556 475 559 524
rect 564 475 567 524
rect 572 475 575 524
rect 580 475 583 524
rect 588 475 591 524
rect 596 475 599 524
rect 604 475 607 524
rect 612 475 615 524
rect 620 475 623 524
rect 628 475 631 524
rect 636 475 639 524
rect 644 475 647 524
rect 652 475 655 524
rect 660 475 663 524
rect 857 518 923 522
rect 927 518 969 522
rect 694 505 735 508
rect 750 505 769 508
rect 672 501 686 502
rect 672 499 724 501
rect 683 498 724 499
rect 732 500 735 505
rect 835 501 871 504
rect 875 501 929 504
rect 933 501 976 504
rect 732 497 769 500
rect 803 492 871 495
rect 875 493 929 496
rect 933 493 976 496
rect 750 489 769 492
rect 672 485 686 486
rect 672 483 724 485
rect 683 482 724 483
rect 835 485 871 488
rect 875 485 929 488
rect 933 485 976 488
rect 444 472 448 475
rect 460 472 464 475
rect 468 472 472 475
rect 484 472 488 475
rect 492 472 496 475
rect 500 472 504 475
rect 508 472 512 475
rect 516 472 520 475
rect 524 472 528 475
rect 532 472 536 475
rect 540 472 544 475
rect 548 472 552 475
rect 556 472 560 475
rect 564 472 568 475
rect 572 472 576 475
rect 580 472 584 475
rect 588 472 592 475
rect 596 472 600 475
rect 604 472 608 475
rect 612 472 616 475
rect 620 472 624 475
rect 628 472 632 475
rect 636 472 640 475
rect 644 472 648 475
rect 652 472 656 475
rect 660 472 664 475
rect 711 473 846 476
rect 1071 475 1074 481
rect 1079 475 1082 481
rect 0 408 3 426
rect 8 396 11 444
rect 16 409 19 426
rect 24 404 27 444
rect 32 404 35 426
rect 40 409 43 444
rect 48 409 51 444
rect 56 404 59 426
rect 64 404 67 444
rect 445 468 448 472
rect 461 468 464 472
rect 469 468 472 472
rect 485 468 488 472
rect 493 468 496 472
rect 501 468 504 472
rect 509 468 512 472
rect 517 468 520 472
rect 525 468 528 472
rect 533 468 536 472
rect 541 468 544 472
rect 549 468 552 472
rect 557 468 560 472
rect 565 468 568 472
rect 573 468 576 472
rect 581 468 584 472
rect 589 468 592 472
rect 597 468 600 472
rect 605 468 608 472
rect 613 468 616 472
rect 621 468 624 472
rect 629 468 632 472
rect 637 468 640 472
rect 645 468 648 472
rect 653 468 656 472
rect 661 468 664 472
rect 674 465 689 468
rect 721 465 731 469
rect 735 465 853 469
rect 250 421 389 424
rect 445 423 448 464
rect 461 423 464 464
rect 250 413 389 416
rect 24 401 28 404
rect 32 401 36 404
rect 56 401 60 404
rect 64 401 68 404
rect 77 401 94 404
rect 113 401 220 404
rect 25 396 28 401
rect 33 396 36 401
rect 57 396 60 401
rect 65 396 68 401
rect 79 393 120 397
rect 124 393 134 397
rect 138 393 227 397
rect 25 364 28 392
rect 33 342 36 392
rect 57 364 60 392
rect 65 342 68 392
rect 90 385 163 389
rect 167 385 197 389
rect 224 385 246 388
rect 262 382 265 403
rect 310 382 313 403
rect 469 387 472 464
rect 485 387 488 464
rect 493 423 496 464
rect 501 387 504 464
rect 509 423 512 464
rect 517 387 520 464
rect 525 423 528 464
rect 533 387 536 464
rect 541 423 544 464
rect 549 387 552 464
rect 557 423 560 464
rect 565 387 568 464
rect 573 423 576 464
rect 581 387 584 464
rect 589 423 592 464
rect 597 387 600 464
rect 605 423 608 464
rect 613 387 616 464
rect 621 423 624 464
rect 629 387 632 464
rect 637 423 640 464
rect 645 387 648 464
rect 653 423 656 464
rect 661 387 664 464
rect 685 457 762 461
rect 766 457 806 461
rect 850 451 877 454
rect 674 443 717 447
rect 885 442 888 475
rect 955 442 958 475
rect 995 442 998 475
rect 1041 442 1044 475
rect 1071 472 1075 475
rect 1079 472 1083 475
rect 1072 468 1075 472
rect 1080 468 1083 472
rect 885 439 897 442
rect 955 439 959 442
rect 995 439 1007 442
rect 1041 439 1045 442
rect 842 399 877 402
rect 262 379 274 382
rect 310 379 322 382
rect 216 351 246 354
rect 33 334 36 338
rect 65 334 68 338
rect 24 331 36 334
rect 56 331 68 334
rect 271 331 274 379
rect -21 325 -1 329
rect 24 317 27 331
rect 56 317 59 331
rect 90 320 246 324
rect 31 309 34 313
rect 63 309 66 313
rect -14 303 -1 306
rect 24 306 34 309
rect 56 306 66 309
rect 286 308 289 371
rect 319 331 322 379
rect 334 308 337 371
rect -21 295 -1 299
rect 24 276 27 306
rect 32 264 35 288
rect 56 268 59 306
rect 79 302 101 305
rect 286 305 297 308
rect 334 305 345 308
rect 64 264 67 288
rect 79 275 94 278
rect 224 275 246 278
rect 262 264 265 289
rect 294 264 297 305
rect 310 264 313 289
rect 342 264 345 305
rect 367 293 371 369
rect 469 365 472 383
rect 501 365 504 383
rect 517 365 520 383
rect 533 365 536 383
rect 549 365 552 383
rect 565 365 568 383
rect 581 365 584 383
rect 597 365 600 383
rect 613 365 616 383
rect 629 365 632 383
rect 645 365 648 383
rect 661 365 664 383
rect 894 367 897 439
rect 460 362 472 365
rect 492 362 504 365
rect 508 362 520 365
rect 524 362 536 365
rect 540 362 552 365
rect 556 362 568 365
rect 572 362 584 365
rect 588 362 600 365
rect 604 362 616 365
rect 620 362 632 365
rect 636 362 648 365
rect 652 362 664 365
rect 415 356 435 360
rect 460 348 463 362
rect 492 348 495 362
rect 508 348 511 362
rect 524 348 527 362
rect 540 348 543 362
rect 556 348 559 362
rect 572 348 575 362
rect 588 348 591 362
rect 604 348 607 362
rect 620 348 623 362
rect 636 348 639 362
rect 652 348 655 362
rect 685 356 877 360
rect 451 340 454 344
rect 467 340 470 344
rect 499 340 502 344
rect 515 340 518 344
rect 531 340 534 344
rect 547 340 550 344
rect 563 340 566 344
rect 579 340 582 344
rect 595 340 598 344
rect 611 340 614 344
rect 627 340 630 344
rect 643 340 646 344
rect 659 340 662 344
rect 422 334 435 337
rect 444 337 454 340
rect 460 337 470 340
rect 492 337 502 340
rect 508 337 518 340
rect 524 337 534 340
rect 540 337 550 340
rect 556 337 566 340
rect 572 337 582 340
rect 588 337 598 340
rect 604 337 614 340
rect 620 337 630 340
rect 636 337 646 340
rect 652 337 662 340
rect 415 326 435 330
rect 444 316 447 337
rect 460 316 463 337
rect 422 302 435 305
rect 444 264 447 312
rect 460 264 463 312
rect 468 289 471 319
rect 492 316 495 337
rect 468 261 471 285
rect 492 265 495 312
rect 500 289 503 319
rect 508 316 511 337
rect 500 261 503 285
rect 508 264 511 312
rect 516 289 519 319
rect 524 316 527 337
rect 516 261 519 285
rect 524 265 527 312
rect 532 289 535 319
rect 540 316 543 337
rect 532 261 535 285
rect 540 265 543 312
rect 548 289 551 319
rect 556 316 559 337
rect 548 261 551 285
rect 556 265 559 312
rect 564 289 567 319
rect 572 316 575 337
rect 564 261 567 285
rect 572 265 575 312
rect 580 289 583 319
rect 588 316 591 337
rect 580 261 583 285
rect 588 265 591 312
rect 596 289 599 319
rect 604 316 607 337
rect 596 261 599 285
rect 604 265 607 312
rect 612 289 615 319
rect 620 316 623 337
rect 612 261 615 285
rect 620 265 623 312
rect 628 289 631 319
rect 636 316 639 337
rect 628 261 631 285
rect 636 265 639 312
rect 644 289 647 319
rect 652 316 655 337
rect 674 333 696 336
rect 644 261 647 285
rect 652 265 655 312
rect 660 289 663 319
rect 918 305 922 429
rect 939 332 942 431
rect 1004 367 1007 439
rect 1025 332 1028 431
rect 1072 423 1075 464
rect 1080 387 1083 464
rect 1080 365 1083 383
rect 1071 362 1083 365
rect 1071 348 1074 362
rect 1078 340 1081 344
rect 1071 337 1081 340
rect 939 329 950 332
rect 1025 329 1036 332
rect 674 301 696 304
rect 660 261 663 285
rect 850 281 877 284
rect 674 272 689 275
rect 885 264 888 301
rect 947 264 950 329
rect 955 264 958 301
rect 995 264 998 301
rect 1033 264 1036 329
rect 1071 316 1074 337
rect 1041 264 1044 301
rect 1071 268 1074 312
rect 1079 292 1082 319
rect 1079 264 1082 288
<< labels >>
rlabel space 69 518 77 524 7 Otop-mid
rlabel space 19 512 39 542 0 top-and
rlabel metal1 82 264 90 264 1 Vdd
rlabel metal1 227 264 235 264 1 GND
rlabel metal2 64 264 67 264 1 <input>
rlabel metal1 262 294 265 294 1 <output>
rlabel metal1 310 294 313 294 1 <output>
rlabel metal2 294 294 297 294 1 <output>
rlabel metal2 342 294 345 294 1 <output>
rlabel metal1 94 264 97 264 1 p2
rlabel metal1 102 264 105 264 1 p2-
rlabel metal1 212 264 215 264 1 p1-
rlabel metal1 220 264 223 264 1 p1
rlabel space -26 425 5 456 1 HGleft-and
rlabel space -26 472 5 480 1 leftu-and
rlabel metal1 885 307 888 307 1 <output>
rlabel metal2 947 307 950 307 1 <output>
rlabel metal1 838 265 841 265 1 p1-
rlabel metal1 846 265 849 265 1 p1
rlabel space 667 584 881 615 1 HG-mid
rlabel space 667 615 881 645 1 midd
rlabel metal2 1033 307 1036 307 1 <output>
rlabel metal1 995 307 998 307 1 <output>
rlabel space 667 705 881 725 1 midu
rlabel space 667 669 881 696 1 top-mid
rlabel space 913 667 937 696 1 VGtop-or
rlabel space 3 409 15 417 0 l1-and
rlabel space 19 409 31 417 0 l0-and
rlabel space 11 417 23 425 0 r1-and
rlabel space 27 417 39 425 0 r0-and
rlabel space 35 409 47 417 0 l.-and
rlabel space 43 417 55 425 0 r.-and
rlabel space 19 464 27 472 0 sp-and
rlabel space 19 425 31 456 0 HGl.-and
rlabel space 35 425 47 456 0 HGl-and
rlabel space 43 425 55 456 1 HGr-and
rlabel space 59 425 71 456 0 HGr.-and
rlabel space 372 409 393 421 0 rightd-or
rlabel space 250 409 262 421 0 d1-or
rlabel space 258 409 270 421 0 d0-or
rlabel space 372 417 393 429 0 rightu-or
rlabel space 306 421 314 429 0 sp-or
rlabel space 250 417 262 429 0 u1-or
rlabel space 258 417 270 429 0 u0-or
rlabel space 250 464 262 476 0 u.-or
rlabel space 250 456 262 468 0 d.-or
rlabel space 889 584 901 615 0 HG-or
rlabel space 913 536 935 548 0 VGd-or
rlabel space 913 560 935 572 0 VGu-or
rlabel space 996 562 1018 574 0 VGu.-or
rlabel space 996 538 1018 550 0 VGd.-or
rlabel space 913 584 935 615 0 HVG-or
rlabel space 959 584 980 615 0 HGright-or
rlabel space -26 464 5 472 3 leftd-and
rlabel space 372 516 393 545 1 ur-or
rlabel space 250 516 262 545 1 topl-or
rlabel space 300 516 312 545 1 topr-or
rlabel space -26 512 5 542 1 ul-and
rlabel space 5 512 7 543 1 Oleft-and
rlabel metal2 468 283 471 283 1 <input>
rlabel metal1 697 262 700 262 1 p2-
rlabel metal1 689 262 692 262 1 p2
rlabel space 455 260 477 481 1 Cbot-and
rlabel space 410 260 441 481 1 ll-and
rlabel space 667 260 881 481 1 bot-mid
rlabel space 1066 260 1088 481 1 bot-and
rlabel space 1025 260 1041 481 1 botr-or
rlabel space 991 260 1015 481 1 botl-or
rlabel space 939 260 955 481 1 Cbotr-or
rlabel space 913 260 935 481 1 VGbot-or
rlabel space 959 260 980 481 1 lr-or
rlabel metal1 677 262 685 262 1 Vdd!
rlabel metal1 853 265 861 265 1 GND!
rlabel space 881 260 905 481 1 Cbotl-or
<< end >>
