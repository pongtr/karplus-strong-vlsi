magic
tech scmos
timestamp 1512638031
<< ntransistor >>
rect 42 -30 44 -26
rect 42 -38 44 -34
rect 58 -30 60 -26
rect 66 -30 68 -26
rect 42 -46 44 -42
rect 50 -46 52 -42
rect 42 -54 44 -50
rect 50 -54 52 -50
rect 66 -38 68 -34
rect 90 -6 92 -2
rect 145 5 149 7
rect 185 5 189 7
rect 106 -6 108 -2
rect 156 -3 160 -1
rect 286 0 296 2
rect 177 -3 181 -1
rect 90 -14 92 -10
rect 98 -14 100 -10
rect 82 -22 84 -18
rect 90 -30 92 -26
rect 82 -38 84 -34
rect 74 -46 76 -42
rect 90 -46 92 -42
rect 145 -11 149 -9
rect 347 -3 351 -1
rect 306 -8 316 -6
rect 185 -11 189 -9
rect 106 -22 108 -18
rect 156 -19 160 -17
rect 355 -11 359 -9
rect 363 -11 367 -9
rect 379 -11 383 -9
rect 286 -16 296 -14
rect 177 -19 181 -17
rect 106 -30 108 -26
rect 145 -27 149 -25
rect 355 -19 359 -17
rect 371 -19 375 -17
rect 387 -19 391 -17
rect 306 -24 316 -22
rect 185 -27 189 -25
rect 106 -38 108 -34
rect 156 -35 160 -33
rect 339 -27 343 -25
rect 286 -32 296 -30
rect 177 -35 181 -33
rect 106 -46 108 -42
rect 339 -35 343 -33
rect 306 -40 316 -38
rect 185 -43 189 -41
rect 90 -54 92 -50
rect 98 -54 100 -50
rect 331 -43 335 -41
rect 286 -48 296 -46
rect 177 -51 181 -49
rect 331 -51 335 -49
rect 40 -87 42 -74
rect 32 -110 34 -97
rect 56 -87 58 -74
rect 48 -110 50 -97
rect 72 -87 74 -74
rect 64 -110 66 -97
rect 88 -87 90 -74
rect 80 -110 82 -97
rect 104 -87 106 -74
rect 344 -84 346 -72
rect 96 -110 98 -97
rect 336 -97 338 -87
rect 360 -84 362 -72
rect 352 -97 354 -87
rect 376 -84 378 -72
rect 368 -97 370 -87
rect 336 -251 338 -239
rect 392 -84 394 -72
rect 384 -97 386 -87
rect 352 -251 354 -239
rect 41 -262 45 -260
rect 57 -262 61 -260
rect 73 -262 77 -260
rect 89 -262 93 -260
rect 105 -262 109 -260
rect 41 -267 45 -265
rect 57 -267 61 -265
rect 73 -267 77 -265
rect 89 -267 93 -265
rect 105 -267 109 -265
rect 344 -266 346 -254
rect 368 -251 370 -239
rect 360 -266 362 -254
rect 384 -251 386 -239
rect 376 -266 378 -254
rect 392 -266 394 -254
<< ptransistor >>
rect 331 21 335 23
rect 339 21 343 23
rect 347 21 351 23
rect 355 21 359 23
rect 363 21 367 23
rect 371 21 375 23
rect 379 21 383 23
rect 387 21 391 23
rect 10 -6 12 -2
rect 10 -14 12 -10
rect 10 -22 12 -18
rect 10 -30 12 -26
rect 10 -38 12 -34
rect 10 -46 12 -42
rect 10 -54 12 -50
rect 129 5 133 7
rect 201 5 205 7
rect 129 -3 133 -1
rect 254 0 274 2
rect 201 -3 205 -1
rect 129 -11 133 -9
rect 224 -8 244 -6
rect 201 -11 205 -9
rect 129 -19 133 -17
rect 254 -16 274 -14
rect 201 -19 205 -17
rect 129 -27 133 -25
rect 224 -24 244 -22
rect 201 -27 205 -25
rect 129 -35 133 -33
rect 254 -32 274 -30
rect 201 -35 205 -33
rect 224 -40 244 -38
rect 201 -43 205 -41
rect 254 -48 274 -46
rect 201 -51 205 -49
rect 32 -147 34 -122
rect 48 -147 50 -122
rect 40 -183 42 -157
rect 64 -147 66 -122
rect 56 -183 58 -157
rect 80 -147 82 -122
rect 72 -183 74 -157
rect 96 -147 98 -122
rect 88 -183 90 -157
rect 336 -133 338 -109
rect 352 -133 354 -109
rect 104 -183 106 -157
rect 41 -201 45 -199
rect 57 -201 61 -199
rect 73 -201 77 -199
rect 89 -201 93 -199
rect 105 -201 109 -199
rect 41 -206 45 -204
rect 57 -206 61 -204
rect 73 -206 77 -204
rect 89 -206 93 -204
rect 105 -206 109 -204
rect 344 -160 346 -136
rect 368 -133 370 -109
rect 344 -201 346 -177
rect 41 -233 45 -231
rect 57 -233 61 -231
rect 73 -233 77 -231
rect 89 -233 93 -231
rect 336 -227 338 -205
rect 105 -233 109 -231
rect 41 -238 45 -236
rect 57 -238 61 -236
rect 73 -238 77 -236
rect 89 -238 93 -236
rect 105 -238 109 -236
rect 360 -160 362 -136
rect 384 -133 386 -109
rect 360 -201 362 -177
rect 352 -227 354 -205
rect 376 -160 378 -136
rect 376 -201 378 -177
rect 368 -227 370 -205
rect 392 -160 394 -136
rect 392 -201 394 -177
rect 384 -227 386 -205
<< ndiffusion >>
rect 37 -26 41 1
rect 37 -30 42 -26
rect 44 -30 45 -26
rect 37 -34 41 -30
rect 37 -38 42 -34
rect 44 -38 45 -34
rect 37 -42 41 -38
rect 53 -26 57 1
rect 69 -26 73 1
rect 53 -30 58 -26
rect 60 -30 61 -26
rect 65 -30 66 -26
rect 68 -30 73 -26
rect 53 -42 57 -30
rect 37 -46 42 -42
rect 44 -46 45 -42
rect 49 -46 50 -42
rect 52 -46 57 -42
rect 37 -50 41 -46
rect 53 -50 57 -46
rect 37 -54 42 -50
rect 44 -54 45 -50
rect 49 -54 50 -50
rect 52 -54 57 -50
rect 37 -57 41 -54
rect 53 -57 57 -54
rect 69 -34 73 -30
rect 65 -38 66 -34
rect 68 -38 73 -34
rect 69 -42 73 -38
rect 85 -2 89 1
rect 85 -6 90 -2
rect 92 -6 93 -2
rect 85 -10 89 -6
rect 101 -2 105 1
rect 145 7 149 8
rect 145 3 149 5
rect 185 7 189 8
rect 185 3 189 5
rect 145 0 160 3
rect 156 -1 160 0
rect 101 -6 106 -2
rect 108 -6 109 -2
rect 177 0 189 3
rect 177 -1 181 0
rect 286 2 296 3
rect 101 -10 105 -6
rect 85 -14 90 -10
rect 92 -14 93 -10
rect 97 -14 98 -10
rect 100 -14 105 -10
rect 85 -18 89 -14
rect 81 -22 82 -18
rect 84 -22 89 -18
rect 85 -26 89 -22
rect 85 -30 90 -26
rect 92 -30 93 -26
rect 85 -34 89 -30
rect 81 -38 82 -34
rect 84 -38 89 -34
rect 69 -46 74 -42
rect 76 -46 77 -42
rect 69 -57 73 -46
rect 85 -42 89 -38
rect 85 -46 90 -42
rect 92 -46 93 -42
rect 85 -50 89 -46
rect 101 -18 105 -14
rect 156 -4 160 -3
rect 177 -4 181 -3
rect 156 -7 159 -4
rect 145 -9 149 -8
rect 145 -13 149 -11
rect 185 -9 189 -8
rect 286 -1 296 0
rect 347 -1 351 0
rect 298 -5 299 -1
rect 303 -5 304 -1
rect 314 -5 316 -1
rect 347 -4 351 -3
rect 306 -6 316 -5
rect 327 -8 396 -4
rect 306 -9 316 -8
rect 355 -9 359 -8
rect 363 -9 367 -8
rect 379 -9 383 -8
rect 185 -13 189 -11
rect 145 -16 160 -13
rect 156 -17 160 -16
rect 101 -22 106 -18
rect 108 -22 109 -18
rect 177 -16 189 -13
rect 177 -17 181 -16
rect 355 -12 359 -11
rect 286 -14 296 -13
rect 363 -12 367 -11
rect 379 -12 383 -11
rect 101 -26 105 -22
rect 101 -30 106 -26
rect 108 -30 109 -26
rect 156 -20 160 -19
rect 177 -20 181 -19
rect 156 -23 159 -20
rect 145 -25 149 -24
rect 101 -34 105 -30
rect 145 -29 149 -27
rect 185 -25 189 -24
rect 286 -17 296 -16
rect 355 -17 359 -16
rect 371 -17 375 -16
rect 387 -17 391 -16
rect 298 -21 299 -17
rect 303 -21 304 -17
rect 314 -21 316 -17
rect 355 -20 359 -19
rect 371 -20 375 -19
rect 387 -20 391 -19
rect 306 -22 316 -21
rect 327 -24 396 -20
rect 306 -25 316 -24
rect 339 -25 343 -24
rect 185 -29 189 -27
rect 145 -32 160 -29
rect 156 -33 160 -32
rect 101 -38 106 -34
rect 108 -38 109 -34
rect 177 -32 189 -29
rect 177 -33 181 -32
rect 339 -28 343 -27
rect 286 -30 296 -29
rect 101 -42 105 -38
rect 101 -46 106 -42
rect 108 -46 109 -42
rect 156 -36 160 -35
rect 177 -36 181 -35
rect 156 -39 159 -36
rect 185 -41 189 -40
rect 286 -33 296 -32
rect 339 -33 343 -32
rect 298 -37 299 -33
rect 303 -37 304 -33
rect 314 -37 316 -33
rect 339 -36 343 -35
rect 306 -38 316 -37
rect 327 -40 396 -36
rect 306 -41 316 -40
rect 331 -41 335 -40
rect 185 -45 189 -43
rect 101 -50 105 -46
rect 85 -54 90 -50
rect 92 -54 93 -50
rect 97 -54 98 -50
rect 100 -54 105 -50
rect 85 -57 89 -54
rect 101 -57 105 -54
rect 177 -48 189 -45
rect 177 -49 181 -48
rect 331 -44 335 -43
rect 286 -46 296 -45
rect 177 -52 181 -51
rect 286 -49 296 -48
rect 331 -49 335 -48
rect 298 -53 299 -49
rect 331 -52 335 -51
rect 327 -56 396 -52
rect 347 -70 351 -69
rect 37 -76 40 -74
rect 39 -87 40 -76
rect 42 -87 43 -74
rect 53 -76 56 -74
rect 35 -90 39 -89
rect 35 -95 39 -94
rect 31 -110 32 -97
rect 34 -110 35 -97
rect 55 -87 56 -76
rect 58 -87 59 -74
rect 69 -76 72 -74
rect 51 -90 55 -89
rect 51 -95 55 -94
rect 47 -110 48 -97
rect 50 -110 51 -97
rect 71 -87 72 -76
rect 74 -87 75 -74
rect 85 -76 88 -74
rect 67 -90 71 -89
rect 67 -95 71 -94
rect 63 -110 64 -97
rect 66 -110 67 -97
rect 87 -87 88 -76
rect 90 -87 91 -74
rect 101 -76 104 -74
rect 83 -90 87 -89
rect 83 -95 87 -94
rect 79 -110 80 -97
rect 82 -110 83 -97
rect 103 -87 104 -76
rect 106 -87 107 -74
rect 340 -84 344 -72
rect 346 -79 347 -72
rect 363 -70 367 -69
rect 346 -84 350 -79
rect 340 -87 343 -84
rect 99 -90 103 -89
rect 99 -95 103 -94
rect 95 -110 96 -97
rect 98 -110 99 -97
rect 332 -89 336 -87
rect 335 -97 336 -89
rect 338 -97 343 -87
rect 356 -84 360 -72
rect 362 -79 363 -72
rect 379 -70 383 -69
rect 362 -84 366 -79
rect 356 -87 359 -84
rect 348 -89 352 -87
rect 351 -97 352 -89
rect 354 -97 359 -87
rect 372 -84 376 -72
rect 378 -79 379 -72
rect 395 -70 399 -69
rect 378 -84 382 -79
rect 372 -87 375 -84
rect 364 -89 368 -87
rect 367 -97 368 -89
rect 370 -97 375 -87
rect 335 -249 336 -239
rect 332 -251 336 -249
rect 338 -251 343 -239
rect 47 -259 48 -255
rect 41 -260 45 -259
rect 63 -259 64 -255
rect 57 -260 61 -259
rect 79 -259 80 -255
rect 73 -260 77 -259
rect 95 -259 96 -255
rect 89 -260 93 -259
rect 111 -259 112 -255
rect 340 -254 343 -251
rect 388 -84 392 -72
rect 394 -79 395 -72
rect 394 -84 398 -79
rect 388 -87 391 -84
rect 380 -89 384 -87
rect 383 -97 384 -89
rect 386 -97 391 -87
rect 351 -249 352 -239
rect 348 -251 352 -249
rect 354 -251 359 -239
rect 105 -260 109 -259
rect 41 -265 45 -262
rect 57 -265 61 -262
rect 73 -265 77 -262
rect 89 -265 93 -262
rect 105 -265 109 -262
rect 41 -268 45 -267
rect 41 -271 42 -268
rect 57 -268 61 -267
rect 57 -271 58 -268
rect 73 -268 77 -267
rect 73 -271 74 -268
rect 89 -268 93 -267
rect 89 -271 90 -268
rect 340 -266 344 -254
rect 346 -259 350 -254
rect 356 -254 359 -251
rect 367 -249 368 -239
rect 364 -251 368 -249
rect 370 -251 375 -239
rect 346 -266 347 -259
rect 105 -268 109 -267
rect 356 -266 360 -254
rect 362 -259 366 -254
rect 372 -254 375 -251
rect 383 -249 384 -239
rect 380 -251 384 -249
rect 386 -251 391 -239
rect 362 -266 363 -259
rect 372 -266 376 -254
rect 378 -259 382 -254
rect 388 -254 391 -251
rect 378 -266 379 -259
rect 388 -266 392 -254
rect 394 -259 398 -254
rect 394 -266 395 -259
rect 105 -271 106 -268
rect 347 -269 351 -268
rect 363 -269 367 -268
rect 379 -269 383 -268
rect 395 -269 399 -268
<< pdiffusion >>
rect 329 28 393 29
rect 331 23 335 24
rect 339 23 343 24
rect 347 23 351 24
rect 355 23 359 24
rect 363 23 367 24
rect 371 23 375 24
rect 379 23 383 24
rect 387 23 391 24
rect 331 20 335 21
rect 339 20 343 21
rect 347 20 351 21
rect 355 20 359 21
rect 363 20 367 21
rect 371 20 375 21
rect 379 20 383 21
rect 387 20 391 21
rect 126 8 127 12
rect 4 -56 5 0
rect 9 -6 10 -2
rect 12 -6 13 -2
rect 9 -14 10 -10
rect 12 -14 13 -10
rect 9 -22 10 -18
rect 12 -22 13 -18
rect 9 -30 10 -26
rect 12 -30 13 -26
rect 9 -38 10 -34
rect 12 -38 13 -34
rect 9 -46 10 -42
rect 12 -46 13 -42
rect 9 -54 10 -50
rect 12 -54 13 -50
rect 129 7 133 8
rect 129 4 133 5
rect 207 8 208 12
rect 201 7 205 8
rect 129 -1 133 0
rect 201 4 205 5
rect 254 3 259 7
rect 201 -1 205 0
rect 254 2 274 3
rect 254 -1 274 0
rect 129 -4 133 -3
rect 201 -4 205 -3
rect 126 -8 127 -4
rect 129 -9 133 -8
rect 129 -12 133 -11
rect 207 -8 208 -4
rect 224 -5 226 -1
rect 246 -5 247 -1
rect 251 -5 252 -1
rect 201 -9 205 -8
rect 224 -6 244 -5
rect 224 -9 244 -8
rect 129 -17 133 -16
rect 201 -12 205 -11
rect 224 -13 226 -9
rect 254 -13 259 -9
rect 201 -17 205 -16
rect 254 -14 274 -13
rect 254 -17 274 -16
rect 129 -20 133 -19
rect 201 -20 205 -19
rect 126 -24 127 -20
rect 129 -25 133 -24
rect 129 -28 133 -27
rect 207 -24 208 -20
rect 224 -21 226 -17
rect 246 -21 247 -17
rect 251 -21 252 -17
rect 201 -25 205 -24
rect 224 -22 244 -21
rect 224 -25 244 -24
rect 129 -33 133 -32
rect 201 -28 205 -27
rect 224 -29 226 -25
rect 254 -29 259 -25
rect 201 -33 205 -32
rect 254 -30 274 -29
rect 254 -33 274 -32
rect 129 -36 133 -35
rect 126 -40 127 -36
rect 201 -36 205 -35
rect 207 -40 208 -36
rect 224 -37 226 -33
rect 246 -37 247 -33
rect 251 -37 252 -33
rect 201 -41 205 -40
rect 224 -38 244 -37
rect 224 -41 244 -40
rect 201 -44 205 -43
rect 224 -45 226 -41
rect 254 -45 259 -41
rect 201 -49 205 -48
rect 254 -46 274 -45
rect 254 -49 274 -48
rect 201 -52 205 -51
rect 207 -56 208 -52
rect 251 -53 252 -49
rect 31 -140 32 -122
rect 29 -147 32 -140
rect 34 -147 35 -122
rect 35 -150 39 -149
rect 35 -155 39 -154
rect 47 -140 48 -122
rect 45 -147 48 -140
rect 50 -147 51 -122
rect 39 -181 40 -157
rect 35 -183 40 -181
rect 42 -174 43 -157
rect 42 -183 45 -174
rect 51 -150 55 -149
rect 51 -155 55 -154
rect 63 -140 64 -122
rect 61 -147 64 -140
rect 66 -147 67 -122
rect 55 -181 56 -157
rect 51 -183 56 -181
rect 58 -174 59 -157
rect 58 -183 61 -174
rect 67 -150 71 -149
rect 67 -155 71 -154
rect 79 -140 80 -122
rect 77 -147 80 -140
rect 82 -147 83 -122
rect 71 -181 72 -157
rect 67 -183 72 -181
rect 74 -174 75 -157
rect 74 -183 77 -174
rect 83 -150 87 -149
rect 83 -155 87 -154
rect 95 -140 96 -122
rect 93 -147 96 -140
rect 98 -147 99 -122
rect 87 -181 88 -157
rect 83 -183 88 -181
rect 90 -174 91 -157
rect 90 -183 93 -174
rect 99 -150 103 -149
rect 99 -155 103 -154
rect 335 -131 336 -109
rect 332 -133 336 -131
rect 338 -133 343 -109
rect 340 -136 343 -133
rect 351 -131 352 -109
rect 348 -133 352 -131
rect 354 -133 359 -109
rect 103 -181 104 -157
rect 99 -183 104 -181
rect 106 -174 107 -157
rect 106 -183 109 -174
rect 41 -198 42 -196
rect 41 -199 45 -198
rect 57 -198 58 -196
rect 57 -199 61 -198
rect 73 -198 74 -196
rect 73 -199 77 -198
rect 89 -198 90 -196
rect 89 -199 93 -198
rect 105 -198 106 -196
rect 105 -199 109 -198
rect 41 -204 45 -201
rect 57 -204 61 -201
rect 73 -204 77 -201
rect 89 -204 93 -201
rect 105 -204 109 -201
rect 340 -160 344 -136
rect 346 -141 350 -136
rect 356 -136 359 -133
rect 367 -131 368 -109
rect 364 -133 368 -131
rect 370 -133 375 -109
rect 346 -160 347 -141
rect 347 -163 351 -162
rect 340 -201 344 -177
rect 346 -201 347 -177
rect 340 -205 343 -201
rect 41 -207 45 -206
rect 47 -211 48 -207
rect 57 -207 61 -206
rect 63 -211 64 -207
rect 73 -207 77 -206
rect 79 -211 80 -207
rect 89 -207 93 -206
rect 95 -211 96 -207
rect 105 -207 109 -206
rect 111 -211 112 -207
rect 41 -230 42 -228
rect 41 -231 45 -230
rect 57 -230 58 -228
rect 57 -231 61 -230
rect 73 -230 74 -228
rect 73 -231 77 -230
rect 89 -230 90 -228
rect 89 -231 93 -230
rect 105 -230 106 -228
rect 335 -227 336 -205
rect 338 -227 343 -205
rect 105 -231 109 -230
rect 41 -236 45 -233
rect 57 -236 61 -233
rect 73 -236 77 -233
rect 89 -236 93 -233
rect 105 -236 109 -233
rect 41 -239 45 -238
rect 47 -243 48 -239
rect 57 -239 61 -238
rect 63 -243 64 -239
rect 73 -239 77 -238
rect 79 -243 80 -239
rect 89 -239 93 -238
rect 95 -243 96 -239
rect 105 -239 109 -238
rect 111 -243 112 -239
rect 356 -160 360 -136
rect 362 -141 366 -136
rect 372 -136 375 -133
rect 383 -131 384 -109
rect 380 -133 384 -131
rect 386 -133 391 -109
rect 362 -160 363 -141
rect 363 -163 367 -162
rect 356 -201 360 -177
rect 362 -201 363 -177
rect 356 -205 359 -201
rect 351 -227 352 -205
rect 354 -227 359 -205
rect 372 -160 376 -136
rect 378 -141 382 -136
rect 388 -136 391 -133
rect 378 -160 379 -141
rect 379 -163 383 -162
rect 372 -201 376 -177
rect 378 -201 379 -177
rect 372 -205 375 -201
rect 367 -227 368 -205
rect 370 -227 375 -205
rect 388 -160 392 -136
rect 394 -141 398 -136
rect 394 -160 395 -141
rect 395 -163 399 -162
rect 388 -201 392 -177
rect 394 -201 395 -177
rect 388 -205 391 -201
rect 383 -227 384 -205
rect 386 -227 391 -205
<< ndcontact >>
rect 37 1 41 5
rect 45 -30 49 -26
rect 45 -38 49 -34
rect 53 1 57 5
rect 69 1 73 5
rect 61 -30 65 -26
rect 45 -46 49 -42
rect 45 -54 49 -50
rect 37 -61 41 -57
rect 53 -61 57 -57
rect 61 -38 65 -34
rect 85 1 89 5
rect 93 -6 97 -2
rect 101 1 105 5
rect 145 8 149 12
rect 185 8 189 12
rect 109 -6 113 -2
rect 286 3 296 7
rect 347 0 351 4
rect 93 -14 97 -10
rect 77 -22 81 -18
rect 93 -30 97 -26
rect 77 -38 81 -34
rect 77 -46 81 -42
rect 69 -61 73 -57
rect 93 -46 97 -42
rect 145 -8 149 -4
rect 159 -8 163 -4
rect 177 -8 181 -4
rect 185 -8 189 -4
rect 286 -5 298 -1
rect 304 -5 314 -1
rect 396 -8 400 -4
rect 109 -22 113 -18
rect 286 -13 296 -9
rect 306 -13 316 -9
rect 355 -16 359 -12
rect 363 -16 367 -12
rect 371 -16 375 -12
rect 379 -16 383 -12
rect 387 -16 391 -12
rect 109 -30 113 -26
rect 145 -24 149 -20
rect 159 -24 163 -20
rect 177 -24 181 -20
rect 185 -24 189 -20
rect 286 -21 298 -17
rect 304 -21 314 -17
rect 396 -24 400 -20
rect 109 -38 113 -34
rect 286 -29 296 -25
rect 306 -29 316 -25
rect 339 -32 343 -28
rect 109 -46 113 -42
rect 159 -40 163 -36
rect 177 -40 181 -36
rect 185 -40 189 -36
rect 286 -37 298 -33
rect 304 -37 314 -33
rect 396 -40 400 -36
rect 93 -54 97 -50
rect 85 -61 89 -57
rect 101 -61 105 -57
rect 286 -45 296 -41
rect 306 -45 316 -41
rect 331 -48 335 -44
rect 177 -56 181 -52
rect 286 -53 298 -49
rect 396 -56 400 -52
rect 35 -89 39 -76
rect 43 -87 47 -74
rect 27 -110 31 -97
rect 35 -110 39 -95
rect 51 -89 55 -76
rect 59 -87 63 -74
rect 43 -110 47 -97
rect 51 -110 55 -95
rect 67 -89 71 -76
rect 75 -87 79 -74
rect 59 -110 63 -97
rect 67 -110 71 -95
rect 83 -89 87 -76
rect 91 -87 95 -74
rect 75 -110 79 -97
rect 83 -110 87 -95
rect 99 -89 103 -76
rect 107 -87 111 -74
rect 347 -79 351 -70
rect 91 -110 95 -97
rect 99 -110 103 -95
rect 331 -97 335 -89
rect 107 -110 111 -97
rect 363 -79 367 -70
rect 347 -97 351 -89
rect 379 -79 383 -70
rect 363 -97 367 -89
rect 331 -249 335 -239
rect 41 -259 47 -255
rect 57 -259 63 -255
rect 73 -259 79 -255
rect 89 -259 95 -255
rect 105 -259 111 -255
rect 395 -79 399 -70
rect 379 -97 383 -89
rect 347 -249 351 -239
rect 42 -272 46 -268
rect 58 -272 62 -268
rect 74 -272 78 -268
rect 90 -272 94 -268
rect 363 -249 367 -239
rect 347 -268 351 -259
rect 379 -249 383 -239
rect 363 -268 367 -259
rect 379 -268 383 -259
rect 395 -268 399 -259
rect 106 -272 110 -268
<< pdcontact >>
rect 329 24 393 28
rect 331 16 335 20
rect 339 16 343 20
rect 347 16 351 20
rect 355 16 359 20
rect 363 16 367 20
rect 371 16 375 20
rect 379 16 383 20
rect 387 16 391 20
rect 127 8 133 12
rect 5 -56 9 0
rect 13 -6 17 -2
rect 13 -14 17 -10
rect 13 -22 17 -18
rect 13 -30 17 -26
rect 13 -38 17 -34
rect 13 -46 17 -42
rect 13 -54 17 -50
rect 129 0 133 4
rect 201 8 207 12
rect 201 0 205 4
rect 259 3 274 7
rect 127 -8 133 -4
rect 129 -16 133 -12
rect 201 -8 207 -4
rect 226 -5 246 -1
rect 252 -5 274 -1
rect 201 -16 205 -12
rect 226 -13 244 -9
rect 259 -13 274 -9
rect 127 -24 133 -20
rect 129 -32 133 -28
rect 201 -24 207 -20
rect 226 -21 246 -17
rect 252 -21 274 -17
rect 201 -32 205 -28
rect 226 -29 244 -25
rect 259 -29 274 -25
rect 127 -40 133 -36
rect 201 -40 207 -36
rect 226 -37 246 -33
rect 252 -37 274 -33
rect 201 -48 205 -44
rect 226 -45 244 -41
rect 259 -45 274 -41
rect 201 -56 207 -52
rect 252 -53 274 -49
rect 27 -140 31 -122
rect 35 -149 39 -122
rect 35 -181 39 -155
rect 43 -140 47 -122
rect 43 -174 47 -155
rect 51 -149 55 -122
rect 51 -181 55 -155
rect 59 -140 63 -122
rect 59 -174 63 -155
rect 67 -149 71 -122
rect 67 -181 71 -155
rect 75 -140 79 -122
rect 75 -174 79 -155
rect 83 -149 87 -122
rect 83 -181 87 -155
rect 91 -140 95 -122
rect 91 -174 95 -155
rect 99 -149 103 -122
rect 99 -181 103 -155
rect 107 -140 111 -122
rect 331 -131 335 -109
rect 347 -131 351 -109
rect 107 -174 111 -155
rect 42 -198 46 -194
rect 58 -198 62 -194
rect 74 -198 78 -194
rect 90 -198 94 -194
rect 106 -198 110 -194
rect 363 -131 367 -109
rect 347 -162 351 -141
rect 347 -201 351 -177
rect 41 -211 47 -207
rect 57 -211 63 -207
rect 73 -211 79 -207
rect 89 -211 95 -207
rect 105 -211 111 -207
rect 42 -230 46 -226
rect 58 -230 62 -226
rect 74 -230 78 -226
rect 90 -230 94 -226
rect 106 -230 110 -226
rect 331 -227 335 -205
rect 41 -243 47 -239
rect 57 -243 63 -239
rect 73 -243 79 -239
rect 89 -243 95 -239
rect 105 -243 111 -239
rect 379 -131 383 -109
rect 363 -162 367 -141
rect 363 -201 367 -177
rect 347 -227 351 -205
rect 379 -162 383 -141
rect 379 -201 383 -177
rect 363 -227 367 -205
rect 395 -162 399 -141
rect 395 -201 399 -177
rect 379 -227 383 -205
<< psubstratepcontact >>
rect 29 26 113 30
rect 396 0 400 4
rect 299 -5 303 -1
rect 396 -16 400 -12
rect 299 -21 303 -17
rect 396 -32 400 -28
rect 299 -37 303 -33
rect 396 -48 400 -44
rect 299 -53 303 -49
rect 299 -64 307 -60
rect 331 -69 335 -65
rect 347 -69 351 -65
rect 35 -94 39 -90
rect 51 -94 55 -90
rect 67 -94 71 -90
rect 83 -94 87 -90
rect 363 -69 367 -65
rect 99 -94 103 -90
rect 379 -69 383 -65
rect 395 -69 399 -65
rect 32 -259 36 -255
rect 48 -259 52 -255
rect 64 -259 68 -255
rect 80 -259 84 -255
rect 96 -259 100 -255
rect 112 -259 116 -255
rect 331 -273 335 -269
rect 347 -273 351 -269
rect 363 -273 367 -269
rect 379 -273 383 -269
rect 395 -273 399 -269
<< nsubstratencontact >>
rect 329 29 393 33
rect 122 8 126 12
rect 0 -56 4 0
rect 208 8 212 12
rect 122 -8 126 -4
rect 208 -8 212 -4
rect 247 -5 251 -1
rect 122 -24 126 -20
rect 208 -24 212 -20
rect 247 -21 251 -17
rect 122 -40 126 -36
rect 208 -40 212 -36
rect 247 -37 251 -33
rect 208 -56 212 -52
rect 247 -53 251 -49
rect 35 -154 39 -150
rect 51 -154 55 -150
rect 67 -154 71 -150
rect 83 -154 87 -150
rect 99 -154 103 -150
rect 331 -167 335 -163
rect 347 -167 351 -163
rect 32 -211 36 -207
rect 48 -211 52 -207
rect 64 -211 68 -207
rect 80 -211 84 -207
rect 96 -211 100 -207
rect 112 -211 116 -207
rect 32 -243 36 -239
rect 48 -243 52 -239
rect 64 -243 68 -239
rect 80 -243 84 -239
rect 96 -243 100 -239
rect 112 -243 116 -239
rect 363 -167 367 -163
rect 379 -167 383 -163
rect 395 -167 399 -163
<< polysilicon >>
rect 324 21 331 23
rect 335 21 339 23
rect 343 21 347 23
rect 351 21 355 23
rect 359 21 363 23
rect 367 21 371 23
rect 375 21 379 23
rect 383 21 387 23
rect 391 21 398 23
rect 10 -2 12 3
rect 10 -10 12 -6
rect 10 -18 12 -14
rect 10 -26 12 -22
rect 10 -34 12 -30
rect 10 -42 12 -38
rect 10 -50 12 -46
rect 10 -59 12 -54
rect 34 -64 36 8
rect 42 -26 44 8
rect 42 -34 44 -30
rect 42 -42 44 -38
rect 50 -42 52 8
rect 58 -26 60 8
rect 66 -26 68 8
rect 42 -50 44 -46
rect 50 -50 52 -46
rect 42 -64 44 -54
rect 50 -64 52 -54
rect 58 -64 60 -30
rect 66 -34 68 -30
rect 66 -64 68 -38
rect 74 -42 76 8
rect 82 -18 84 8
rect 90 -2 92 8
rect 90 -10 92 -6
rect 98 -10 100 8
rect 106 -2 108 8
rect 127 5 129 7
rect 133 5 145 7
rect 149 5 152 7
rect 156 5 185 7
rect 189 5 201 7
rect 205 5 207 7
rect 119 -3 129 -1
rect 133 -3 156 -1
rect 160 -3 162 -1
rect 223 0 254 2
rect 274 0 286 2
rect 296 0 298 2
rect 174 -3 177 -1
rect 181 -3 201 -1
rect 205 -3 207 -1
rect 82 -34 84 -22
rect 90 -26 92 -14
rect 74 -64 76 -46
rect 82 -64 84 -38
rect 90 -42 92 -30
rect 90 -50 92 -46
rect 98 -50 100 -14
rect 106 -18 108 -6
rect 119 -12 121 -3
rect 127 -11 129 -9
rect 133 -11 145 -9
rect 149 -11 152 -9
rect 326 -3 347 -1
rect 351 -3 403 -1
rect 223 -8 224 -6
rect 244 -8 306 -6
rect 316 -8 318 -6
rect 156 -11 185 -9
rect 189 -11 201 -9
rect 205 -11 207 -9
rect 119 -19 129 -17
rect 133 -19 156 -17
rect 160 -19 162 -17
rect 326 -11 355 -9
rect 359 -11 363 -9
rect 367 -11 379 -9
rect 383 -11 403 -9
rect 223 -16 254 -14
rect 274 -16 286 -14
rect 296 -16 298 -14
rect 174 -19 177 -17
rect 181 -19 201 -17
rect 205 -19 207 -17
rect 106 -26 108 -22
rect 119 -28 121 -19
rect 127 -27 129 -25
rect 133 -27 145 -25
rect 149 -27 152 -25
rect 106 -34 108 -30
rect 326 -19 355 -17
rect 359 -19 371 -17
rect 375 -19 387 -17
rect 391 -19 403 -17
rect 223 -24 224 -22
rect 244 -24 306 -22
rect 316 -24 318 -22
rect 156 -27 185 -25
rect 189 -27 201 -25
rect 205 -27 207 -25
rect 119 -35 129 -33
rect 133 -35 156 -33
rect 160 -35 162 -33
rect 326 -27 339 -25
rect 343 -27 403 -25
rect 223 -32 254 -30
rect 274 -32 286 -30
rect 296 -32 298 -30
rect 174 -35 177 -33
rect 181 -35 201 -33
rect 205 -35 207 -33
rect 106 -42 108 -38
rect 119 -44 121 -35
rect 326 -35 339 -33
rect 343 -35 403 -33
rect 223 -40 224 -38
rect 244 -40 306 -38
rect 316 -40 318 -38
rect 156 -43 185 -41
rect 189 -43 201 -41
rect 205 -43 207 -41
rect 90 -64 92 -54
rect 98 -64 100 -54
rect 106 -64 108 -46
rect 326 -43 331 -41
rect 335 -43 403 -41
rect 223 -48 254 -46
rect 274 -48 286 -46
rect 296 -48 298 -46
rect 174 -51 177 -49
rect 181 -51 201 -49
rect 205 -51 207 -49
rect 326 -51 331 -49
rect 335 -51 403 -49
rect 343 -62 346 -60
rect 359 -62 362 -60
rect 375 -62 378 -60
rect 391 -62 394 -60
rect 344 -72 346 -62
rect 40 -74 42 -72
rect 56 -74 58 -72
rect 72 -74 74 -72
rect 88 -74 90 -72
rect 104 -74 106 -72
rect 32 -97 34 -95
rect 32 -122 34 -110
rect 32 -184 34 -147
rect 40 -157 42 -87
rect 48 -97 50 -95
rect 48 -122 50 -110
rect 40 -184 42 -183
rect 48 -184 50 -147
rect 56 -157 58 -87
rect 64 -97 66 -95
rect 64 -122 66 -110
rect 56 -184 58 -183
rect 64 -184 66 -147
rect 72 -157 74 -87
rect 80 -97 82 -95
rect 80 -122 82 -110
rect 72 -184 74 -183
rect 80 -184 82 -147
rect 88 -157 90 -87
rect 360 -72 362 -62
rect 336 -87 338 -86
rect 96 -97 98 -95
rect 96 -122 98 -110
rect 88 -184 90 -183
rect 96 -184 98 -147
rect 104 -157 106 -87
rect 336 -101 338 -97
rect 336 -109 338 -107
rect 336 -134 338 -133
rect 344 -136 346 -84
rect 376 -72 378 -62
rect 352 -87 354 -86
rect 352 -101 354 -97
rect 352 -109 354 -107
rect 352 -134 354 -133
rect 104 -184 106 -183
rect 39 -200 41 -199
rect 36 -201 41 -200
rect 45 -201 47 -199
rect 55 -200 57 -199
rect 52 -201 57 -200
rect 61 -201 63 -199
rect 71 -200 73 -199
rect 68 -201 73 -200
rect 77 -201 79 -199
rect 87 -200 89 -199
rect 84 -201 89 -200
rect 93 -201 95 -199
rect 103 -200 105 -199
rect 100 -201 105 -200
rect 109 -201 111 -199
rect 38 -206 41 -204
rect 45 -206 47 -204
rect 54 -206 57 -204
rect 61 -206 63 -204
rect 70 -206 73 -204
rect 77 -206 79 -204
rect 86 -206 89 -204
rect 93 -206 95 -204
rect 102 -206 105 -204
rect 109 -206 111 -204
rect 336 -205 338 -138
rect 360 -136 362 -84
rect 392 -72 394 -62
rect 368 -87 370 -86
rect 368 -101 370 -97
rect 368 -109 370 -107
rect 368 -134 370 -133
rect 344 -162 346 -160
rect 344 -177 346 -174
rect 38 -214 40 -206
rect 54 -214 56 -206
rect 70 -214 72 -206
rect 86 -214 88 -206
rect 102 -214 104 -206
rect 39 -232 41 -231
rect 36 -233 41 -232
rect 45 -233 47 -231
rect 55 -232 57 -231
rect 52 -233 57 -232
rect 61 -233 63 -231
rect 71 -232 73 -231
rect 68 -233 73 -232
rect 77 -233 79 -231
rect 87 -232 89 -231
rect 84 -233 89 -232
rect 93 -233 95 -231
rect 336 -231 338 -227
rect 103 -232 105 -231
rect 100 -233 105 -232
rect 109 -233 111 -231
rect 38 -238 41 -236
rect 45 -238 47 -236
rect 54 -238 57 -236
rect 61 -238 63 -236
rect 70 -238 73 -236
rect 77 -238 79 -236
rect 86 -238 89 -236
rect 93 -238 95 -236
rect 102 -238 105 -236
rect 109 -238 111 -236
rect 38 -248 40 -238
rect 54 -248 56 -238
rect 70 -248 72 -238
rect 86 -248 88 -238
rect 102 -248 104 -238
rect 336 -239 338 -237
rect 336 -252 338 -251
rect 38 -260 40 -252
rect 54 -260 56 -252
rect 70 -260 72 -252
rect 86 -260 88 -252
rect 102 -260 104 -252
rect 344 -254 346 -201
rect 352 -205 354 -138
rect 376 -136 378 -84
rect 384 -87 386 -86
rect 384 -101 386 -97
rect 384 -109 386 -107
rect 384 -134 386 -133
rect 360 -162 362 -160
rect 360 -177 362 -174
rect 352 -231 354 -227
rect 352 -239 354 -237
rect 352 -252 354 -251
rect 38 -262 41 -260
rect 45 -262 47 -260
rect 54 -262 57 -260
rect 61 -262 63 -260
rect 70 -262 73 -260
rect 77 -262 79 -260
rect 86 -262 89 -260
rect 93 -262 95 -260
rect 102 -262 105 -260
rect 109 -262 111 -260
rect 37 -266 41 -265
rect 39 -267 41 -266
rect 45 -267 47 -265
rect 53 -266 57 -265
rect 55 -267 57 -266
rect 61 -267 63 -265
rect 69 -266 73 -265
rect 71 -267 73 -266
rect 77 -267 79 -265
rect 85 -266 89 -265
rect 87 -267 89 -266
rect 93 -267 95 -265
rect 101 -266 105 -265
rect 103 -267 105 -266
rect 109 -267 111 -265
rect 360 -254 362 -201
rect 368 -205 370 -138
rect 392 -136 394 -84
rect 376 -162 378 -160
rect 376 -177 378 -174
rect 368 -231 370 -227
rect 368 -239 370 -237
rect 368 -252 370 -251
rect 344 -268 346 -266
rect 376 -254 378 -201
rect 384 -205 386 -138
rect 392 -162 394 -160
rect 392 -177 394 -174
rect 384 -231 386 -227
rect 384 -239 386 -237
rect 384 -252 386 -251
rect 360 -268 362 -266
rect 392 -254 394 -201
rect 376 -268 378 -266
rect 392 -268 394 -266
<< polycontact >>
rect 398 21 402 25
rect 322 17 326 21
rect 34 8 38 12
rect 42 8 46 12
rect 50 8 54 12
rect 58 8 62 12
rect 66 8 70 12
rect 74 8 78 12
rect 82 8 86 12
rect 90 8 94 12
rect 98 8 102 12
rect 106 8 110 12
rect 8 3 12 7
rect 8 -63 12 -59
rect 152 4 156 8
rect 170 -3 174 1
rect 219 -1 223 3
rect 115 -13 119 -9
rect 152 -12 156 -8
rect 322 -5 326 -1
rect 219 -9 223 -5
rect 403 -5 407 -1
rect 170 -19 174 -15
rect 219 -17 223 -13
rect 322 -13 326 -9
rect 403 -13 407 -9
rect 115 -29 119 -25
rect 152 -28 156 -24
rect 322 -21 326 -17
rect 219 -25 223 -21
rect 403 -21 407 -17
rect 170 -35 174 -31
rect 219 -33 223 -29
rect 322 -29 326 -25
rect 403 -29 407 -25
rect 115 -45 119 -41
rect 152 -44 156 -40
rect 322 -37 326 -33
rect 219 -41 223 -37
rect 403 -37 407 -33
rect 170 -51 174 -47
rect 219 -49 223 -45
rect 322 -45 326 -41
rect 403 -45 407 -41
rect 322 -53 326 -49
rect 403 -53 407 -49
rect 339 -62 343 -58
rect 355 -62 359 -58
rect 371 -62 375 -58
rect 387 -62 391 -58
rect 34 -68 38 -64
rect 42 -68 46 -64
rect 50 -68 54 -64
rect 58 -68 62 -64
rect 66 -68 70 -64
rect 74 -68 78 -64
rect 82 -68 86 -64
rect 90 -68 94 -64
rect 98 -68 102 -64
rect 106 -68 110 -64
rect 335 -86 339 -82
rect 335 -138 339 -134
rect 351 -86 355 -82
rect 32 -188 36 -184
rect 40 -188 44 -184
rect 48 -188 52 -184
rect 56 -188 60 -184
rect 64 -188 68 -184
rect 72 -188 76 -184
rect 80 -188 84 -184
rect 88 -188 92 -184
rect 96 -188 100 -184
rect 104 -188 108 -184
rect 35 -200 39 -196
rect 51 -200 55 -196
rect 67 -200 71 -196
rect 83 -200 87 -196
rect 99 -200 103 -196
rect 351 -138 355 -134
rect 367 -86 371 -82
rect 344 -174 348 -170
rect 37 -218 41 -214
rect 53 -218 57 -214
rect 69 -218 73 -214
rect 85 -218 89 -214
rect 101 -218 105 -214
rect 35 -232 39 -228
rect 51 -232 55 -228
rect 67 -232 71 -228
rect 83 -232 87 -228
rect 99 -232 103 -228
rect 37 -252 41 -248
rect 53 -252 57 -248
rect 69 -252 73 -248
rect 85 -252 89 -248
rect 101 -252 105 -248
rect 335 -256 339 -252
rect 367 -138 371 -134
rect 383 -86 387 -82
rect 360 -174 364 -170
rect 35 -270 39 -266
rect 51 -270 55 -266
rect 67 -270 71 -266
rect 83 -270 87 -266
rect 99 -270 103 -266
rect 351 -256 355 -252
rect 383 -138 387 -134
rect 376 -174 380 -170
rect 367 -256 371 -252
rect 392 -174 396 -170
rect 383 -256 387 -252
<< metal1 >>
rect 16 26 29 30
rect 113 26 303 32
rect 329 28 393 29
rect 16 24 113 26
rect 16 16 20 24
rect 126 8 127 12
rect 137 8 145 11
rect 153 8 156 12
rect 8 7 12 8
rect 30 2 37 5
rect 41 2 53 5
rect 57 2 69 5
rect 73 2 85 5
rect 89 2 101 5
rect 105 2 109 5
rect 4 -56 5 0
rect 17 -6 93 -3
rect 97 -6 109 -3
rect 113 -6 114 -2
rect 122 -4 126 8
rect 137 4 140 8
rect 133 1 136 4
rect 126 -8 127 -4
rect 137 -8 145 -5
rect 153 -8 156 4
rect 17 -14 93 -11
rect 113 -11 115 -10
rect 97 -13 115 -11
rect 97 -14 116 -13
rect 17 -22 77 -19
rect 81 -22 109 -19
rect 113 -22 114 -18
rect 122 -20 126 -8
rect 137 -12 140 -8
rect 133 -15 136 -12
rect 126 -24 127 -20
rect 137 -24 145 -21
rect 153 -24 156 -12
rect 17 -30 45 -27
rect 49 -30 61 -27
rect 65 -30 93 -27
rect 97 -30 109 -27
rect 113 -29 115 -26
rect 113 -30 116 -29
rect 17 -38 45 -35
rect 49 -38 61 -35
rect 65 -38 77 -35
rect 81 -38 109 -35
rect 113 -38 114 -34
rect 122 -36 126 -24
rect 137 -28 140 -24
rect 133 -31 136 -28
rect 126 -40 127 -36
rect 153 -40 156 -28
rect 17 -46 45 -43
rect 49 -46 77 -43
rect 81 -46 93 -43
rect 97 -46 109 -43
rect 113 -45 115 -42
rect 113 -46 116 -45
rect 17 -54 45 -51
rect 49 -54 93 -51
rect 113 -51 114 -50
rect 97 -54 114 -51
rect 122 -56 126 -40
rect 1 -177 5 -56
rect 30 -61 37 -58
rect 41 -61 53 -58
rect 57 -61 69 -58
rect 73 -61 85 -58
rect 89 -61 101 -58
rect 105 -61 119 -58
rect 122 -60 131 -56
rect 8 -64 12 -63
rect 116 -68 119 -61
rect 1 -207 5 -181
rect 9 -199 12 -68
rect 35 -69 39 -68
rect 43 -69 47 -68
rect 51 -69 55 -68
rect 59 -69 63 -68
rect 67 -69 71 -68
rect 75 -69 79 -68
rect 83 -69 87 -68
rect 91 -69 95 -68
rect 99 -69 103 -68
rect 107 -69 111 -68
rect 43 -74 47 -73
rect 59 -74 63 -73
rect 35 -90 39 -89
rect 75 -74 79 -73
rect 51 -90 55 -89
rect 91 -74 95 -73
rect 67 -90 71 -89
rect 107 -74 111 -73
rect 83 -90 87 -89
rect 123 -76 131 -60
rect 153 -60 156 -44
rect 163 -68 167 26
rect 170 -4 174 -3
rect 177 -4 181 26
rect 208 15 292 19
rect 208 12 212 15
rect 189 8 195 11
rect 207 8 208 12
rect 192 4 195 8
rect 196 1 201 4
rect 208 -4 212 8
rect 252 -1 256 15
rect 299 10 303 26
rect 326 24 329 28
rect 393 24 395 28
rect 318 17 322 20
rect 398 20 402 21
rect 274 4 286 7
rect 277 -1 280 4
rect 299 6 322 10
rect 299 -1 303 6
rect 189 -8 195 -5
rect 207 -8 208 -4
rect 246 -5 247 -1
rect 251 -5 252 -1
rect 298 -5 299 -1
rect 303 -5 304 -1
rect 321 -5 322 -1
rect 170 -20 174 -19
rect 177 -20 181 -8
rect 192 -12 195 -8
rect 196 -15 201 -12
rect 208 -20 212 -8
rect 244 -13 245 -9
rect 252 -17 256 -5
rect 274 -12 286 -9
rect 277 -17 280 -12
rect 299 -17 303 -5
rect 316 -13 317 -9
rect 321 -13 322 -9
rect 189 -24 195 -21
rect 207 -24 208 -20
rect 246 -21 247 -17
rect 251 -21 252 -17
rect 298 -21 299 -17
rect 303 -21 304 -17
rect 321 -21 322 -17
rect 170 -36 174 -35
rect 177 -36 181 -24
rect 192 -28 195 -24
rect 196 -31 201 -28
rect 208 -36 212 -24
rect 244 -29 245 -25
rect 252 -33 256 -21
rect 274 -28 286 -25
rect 277 -33 280 -28
rect 299 -33 303 -21
rect 316 -29 317 -25
rect 321 -29 322 -25
rect 189 -40 195 -37
rect 207 -40 208 -36
rect 246 -37 247 -33
rect 251 -37 252 -33
rect 298 -37 299 -33
rect 303 -37 304 -33
rect 321 -37 322 -33
rect 170 -52 174 -51
rect 177 -52 181 -40
rect 192 -44 195 -40
rect 196 -47 201 -44
rect 208 -52 212 -40
rect 244 -45 245 -41
rect 252 -49 256 -37
rect 274 -44 286 -41
rect 277 -49 280 -44
rect 299 -49 303 -37
rect 316 -45 317 -41
rect 321 -45 322 -41
rect 331 -44 334 16
rect 339 -28 342 16
rect 347 4 350 16
rect 207 -56 208 -52
rect 251 -53 252 -49
rect 298 -53 299 -49
rect 321 -53 322 -49
rect 123 -80 127 -76
rect 99 -90 103 -89
rect 9 -231 12 -203
rect 20 -94 35 -90
rect 39 -94 51 -90
rect 55 -94 67 -90
rect 71 -94 83 -90
rect 87 -94 99 -90
rect 103 -94 116 -90
rect 16 -255 20 -94
rect 35 -95 39 -94
rect 51 -95 55 -94
rect 67 -95 71 -94
rect 83 -95 87 -94
rect 99 -95 103 -94
rect 27 -115 30 -110
rect 27 -118 35 -115
rect 43 -115 46 -110
rect 43 -118 51 -115
rect 59 -115 62 -110
rect 59 -118 67 -115
rect 75 -115 78 -110
rect 75 -118 83 -115
rect 91 -115 94 -110
rect 91 -118 99 -115
rect 27 -122 30 -118
rect 43 -122 46 -118
rect 59 -122 62 -118
rect 75 -122 78 -118
rect 91 -122 94 -118
rect 107 -122 110 -110
rect 29 -147 35 -143
rect 39 -147 51 -143
rect 35 -150 39 -149
rect 55 -147 67 -143
rect 51 -150 55 -149
rect 71 -147 83 -143
rect 67 -150 71 -149
rect 87 -147 99 -143
rect 83 -150 87 -149
rect 123 -143 131 -80
rect 103 -147 131 -143
rect 99 -150 103 -149
rect 35 -155 39 -154
rect 29 -181 35 -177
rect 43 -155 47 -154
rect 51 -155 55 -154
rect 39 -181 51 -177
rect 59 -155 63 -154
rect 67 -155 71 -154
rect 55 -181 67 -177
rect 75 -155 79 -154
rect 83 -155 87 -154
rect 71 -181 83 -177
rect 91 -155 95 -154
rect 99 -155 103 -154
rect 87 -181 99 -177
rect 107 -155 111 -154
rect 123 -177 131 -147
rect 103 -181 127 -177
rect 33 -189 37 -188
rect 41 -189 45 -188
rect 49 -189 53 -188
rect 57 -189 61 -188
rect 65 -189 69 -188
rect 73 -189 77 -188
rect 81 -189 85 -188
rect 89 -189 93 -188
rect 97 -189 101 -188
rect 105 -189 109 -188
rect 42 -194 45 -193
rect 58 -194 61 -193
rect 74 -194 77 -193
rect 90 -194 93 -193
rect 106 -194 109 -193
rect 35 -201 39 -200
rect 51 -201 55 -200
rect 67 -201 71 -200
rect 83 -201 87 -200
rect 99 -201 103 -200
rect 29 -203 116 -201
rect 26 -204 116 -203
rect 123 -207 131 -181
rect 29 -211 32 -207
rect 36 -211 41 -207
rect 47 -211 48 -207
rect 52 -211 57 -207
rect 63 -211 64 -207
rect 68 -211 73 -207
rect 79 -211 80 -207
rect 84 -211 89 -207
rect 95 -211 96 -207
rect 100 -211 105 -207
rect 111 -211 112 -207
rect 116 -211 131 -207
rect 41 -218 42 -214
rect 57 -218 58 -214
rect 73 -218 74 -214
rect 89 -218 90 -214
rect 105 -218 106 -214
rect 38 -225 45 -222
rect 54 -225 61 -222
rect 70 -225 77 -222
rect 86 -225 93 -222
rect 102 -225 109 -222
rect 42 -226 45 -225
rect 58 -226 61 -225
rect 74 -226 77 -225
rect 90 -226 93 -225
rect 106 -226 109 -225
rect 35 -233 39 -232
rect 51 -233 55 -232
rect 67 -233 71 -232
rect 83 -233 87 -232
rect 99 -233 103 -232
rect 29 -235 116 -233
rect 26 -236 116 -235
rect 123 -239 131 -211
rect 29 -243 32 -239
rect 36 -243 41 -239
rect 47 -243 48 -239
rect 52 -243 57 -239
rect 63 -243 64 -239
rect 68 -243 73 -239
rect 79 -243 80 -239
rect 84 -243 89 -239
rect 95 -243 96 -239
rect 100 -243 105 -239
rect 111 -243 112 -239
rect 116 -243 131 -239
rect 41 -252 42 -248
rect 57 -252 58 -248
rect 73 -252 74 -248
rect 89 -252 90 -248
rect 105 -252 106 -248
rect 16 -259 32 -255
rect 36 -259 41 -255
rect 47 -259 48 -255
rect 52 -259 57 -255
rect 63 -259 64 -255
rect 68 -259 73 -255
rect 79 -259 80 -255
rect 84 -259 89 -255
rect 95 -259 96 -255
rect 100 -259 105 -255
rect 111 -259 112 -255
rect 29 -265 116 -262
rect 35 -266 39 -265
rect 51 -266 55 -265
rect 67 -266 71 -265
rect 83 -266 87 -265
rect 99 -266 103 -265
rect 42 -273 45 -272
rect 58 -273 61 -272
rect 74 -273 77 -272
rect 90 -273 93 -272
rect 106 -273 109 -272
rect 38 -276 45 -273
rect 54 -276 61 -273
rect 70 -276 77 -273
rect 86 -276 93 -273
rect 102 -276 109 -273
rect 123 -276 131 -243
rect 177 -68 181 -56
rect 135 -262 138 -72
rect 163 -90 167 -72
rect 208 -76 212 -56
rect 252 -76 256 -53
rect 299 -56 303 -53
rect 331 -56 334 -48
rect 339 -56 342 -32
rect 347 -56 350 0
rect 355 -12 358 16
rect 363 -12 366 16
rect 371 -12 374 16
rect 379 -12 382 16
rect 387 -12 390 16
rect 396 4 400 6
rect 396 -4 400 0
rect 407 -5 408 -1
rect 396 -12 400 -8
rect 407 -13 408 -9
rect 355 -56 358 -16
rect 363 -56 366 -16
rect 371 -56 374 -16
rect 379 -56 382 -16
rect 387 -56 390 -16
rect 396 -20 400 -16
rect 407 -21 408 -17
rect 396 -28 400 -24
rect 407 -29 408 -25
rect 396 -36 400 -32
rect 407 -37 408 -33
rect 396 -44 400 -40
rect 407 -45 408 -41
rect 396 -52 400 -48
rect 407 -53 408 -49
rect 299 -60 307 -56
rect 331 -58 335 -56
rect 339 -58 343 -56
rect 347 -58 351 -56
rect 355 -58 359 -56
rect 363 -58 367 -56
rect 371 -58 375 -56
rect 379 -58 383 -56
rect 387 -58 391 -56
rect 292 -82 295 -64
rect 299 -65 307 -64
rect 299 -68 331 -65
rect 303 -69 331 -68
rect 335 -69 347 -65
rect 351 -69 363 -65
rect 367 -69 379 -65
rect 383 -69 395 -65
rect 303 -72 307 -69
rect 143 -232 146 -204
rect 135 -276 138 -266
rect 143 -276 146 -236
rect 284 -273 287 -138
rect 292 -253 295 -86
rect 292 -273 295 -257
rect 299 -269 307 -72
rect 347 -70 351 -69
rect 363 -70 367 -69
rect 379 -70 383 -69
rect 395 -70 399 -69
rect 327 -86 335 -83
rect 339 -86 351 -83
rect 355 -86 367 -83
rect 371 -86 383 -83
rect 387 -86 399 -83
rect 331 -102 334 -97
rect 347 -102 350 -97
rect 363 -102 366 -97
rect 379 -102 382 -97
rect 331 -109 334 -106
rect 347 -109 350 -106
rect 363 -109 366 -106
rect 379 -109 382 -106
rect 327 -138 335 -135
rect 339 -138 351 -135
rect 355 -138 367 -135
rect 371 -138 383 -135
rect 387 -138 399 -135
rect 347 -163 351 -162
rect 363 -163 367 -162
rect 379 -163 383 -162
rect 395 -163 399 -162
rect 323 -167 331 -163
rect 335 -167 347 -163
rect 351 -167 363 -163
rect 367 -167 379 -163
rect 383 -167 395 -163
rect 323 -177 327 -167
rect 343 -174 344 -170
rect 359 -174 360 -170
rect 375 -174 376 -170
rect 391 -174 392 -170
rect 327 -181 347 -177
rect 351 -181 363 -177
rect 367 -181 379 -177
rect 383 -181 395 -177
rect 331 -232 334 -227
rect 347 -232 350 -227
rect 363 -232 366 -227
rect 379 -232 382 -227
rect 331 -239 334 -236
rect 347 -239 350 -236
rect 363 -239 366 -236
rect 379 -239 382 -236
rect 327 -256 335 -253
rect 339 -256 351 -253
rect 355 -256 367 -253
rect 371 -256 383 -253
rect 387 -256 399 -253
rect 347 -269 351 -268
rect 363 -269 367 -268
rect 379 -269 383 -268
rect 395 -269 399 -268
rect 299 -273 331 -269
rect 335 -273 347 -269
rect 351 -273 363 -269
rect 367 -273 379 -269
rect 383 -273 395 -269
<< m2contact >>
rect 16 12 20 16
rect 34 12 38 16
rect 8 8 12 12
rect 42 12 46 16
rect 50 12 54 16
rect 58 12 62 16
rect 66 12 70 16
rect 74 12 78 16
rect 82 12 86 16
rect 90 12 94 16
rect 98 12 102 16
rect 106 12 110 16
rect 26 1 30 5
rect 114 -6 118 -2
rect 136 0 140 4
rect 114 -22 118 -18
rect 136 -16 140 -12
rect 114 -38 118 -34
rect 136 -32 140 -28
rect 114 -54 118 -50
rect 26 -61 30 -57
rect 8 -68 12 -64
rect 1 -181 5 -177
rect 35 -73 39 -69
rect 43 -73 47 -69
rect 51 -73 55 -69
rect 59 -73 63 -69
rect 67 -73 71 -69
rect 75 -73 79 -69
rect 83 -73 87 -69
rect 91 -73 95 -69
rect 99 -73 103 -69
rect 107 -73 111 -69
rect 116 -72 120 -68
rect 153 -64 157 -60
rect 170 -8 174 -4
rect 292 15 296 19
rect 192 0 196 4
rect 215 -1 219 3
rect 322 24 326 28
rect 314 16 318 20
rect 398 16 402 20
rect 322 6 326 10
rect 277 -5 281 -1
rect 317 -5 321 -1
rect 170 -24 174 -20
rect 192 -16 196 -12
rect 215 -9 219 -5
rect 245 -13 249 -9
rect 215 -17 219 -13
rect 317 -13 321 -9
rect 277 -21 281 -17
rect 317 -21 321 -17
rect 170 -40 174 -36
rect 192 -32 196 -28
rect 215 -25 219 -21
rect 245 -29 249 -25
rect 215 -33 219 -29
rect 317 -29 321 -25
rect 277 -37 281 -33
rect 317 -37 321 -33
rect 170 -56 174 -52
rect 192 -48 196 -44
rect 215 -41 219 -37
rect 245 -45 249 -41
rect 215 -49 219 -45
rect 317 -45 321 -41
rect 277 -53 281 -49
rect 317 -53 321 -49
rect 127 -80 131 -76
rect 8 -203 12 -199
rect 1 -211 5 -207
rect 8 -235 12 -231
rect 16 -94 20 -90
rect 116 -94 120 -90
rect 35 -118 39 -114
rect 51 -118 55 -114
rect 67 -118 71 -114
rect 83 -118 87 -114
rect 99 -118 103 -114
rect 25 -181 29 -177
rect 43 -154 47 -150
rect 59 -154 63 -150
rect 75 -154 79 -150
rect 91 -154 95 -150
rect 107 -154 111 -150
rect 127 -181 131 -177
rect 33 -193 37 -189
rect 41 -193 45 -189
rect 49 -193 53 -189
rect 57 -193 61 -189
rect 65 -193 69 -189
rect 73 -193 77 -189
rect 81 -193 85 -189
rect 89 -193 93 -189
rect 97 -193 101 -189
rect 105 -193 109 -189
rect 25 -203 29 -199
rect 116 -204 120 -200
rect 25 -211 29 -207
rect 42 -218 46 -214
rect 58 -218 62 -214
rect 74 -218 78 -214
rect 90 -218 94 -214
rect 106 -218 110 -214
rect 34 -225 38 -221
rect 50 -225 54 -221
rect 66 -225 70 -221
rect 82 -225 86 -221
rect 98 -225 102 -221
rect 25 -235 29 -231
rect 116 -236 120 -232
rect 42 -252 46 -248
rect 58 -252 62 -248
rect 74 -252 78 -248
rect 90 -252 94 -248
rect 106 -252 110 -248
rect 116 -266 120 -262
rect 34 -277 38 -273
rect 50 -277 54 -273
rect 66 -277 70 -273
rect 82 -277 86 -273
rect 98 -277 102 -273
rect 135 -72 139 -68
rect 163 -72 167 -68
rect 177 -72 181 -68
rect 208 -80 212 -76
rect 396 6 400 10
rect 408 -5 412 -1
rect 408 -13 412 -9
rect 408 -21 412 -17
rect 408 -29 412 -25
rect 408 -37 412 -33
rect 408 -45 412 -41
rect 408 -53 412 -49
rect 252 -80 256 -76
rect 292 -64 296 -60
rect 331 -62 335 -58
rect 347 -62 351 -58
rect 363 -62 367 -58
rect 379 -62 383 -58
rect 163 -94 167 -90
rect 299 -72 303 -68
rect 292 -86 296 -82
rect 284 -138 288 -134
rect 142 -204 146 -200
rect 142 -236 146 -232
rect 135 -266 139 -262
rect 292 -257 296 -253
rect 323 -86 327 -82
rect 331 -106 335 -102
rect 347 -106 351 -102
rect 363 -106 367 -102
rect 379 -106 383 -102
rect 323 -138 327 -134
rect 339 -174 343 -170
rect 355 -174 359 -170
rect 371 -174 375 -170
rect 387 -174 391 -170
rect 323 -181 327 -177
rect 331 -236 335 -232
rect 347 -236 351 -232
rect 363 -236 367 -232
rect 379 -236 383 -232
rect 323 -257 327 -253
<< metal2 >>
rect 113 23 280 25
rect 9 22 280 23
rect 9 20 117 22
rect 9 12 12 20
rect 9 -64 12 8
rect 16 -90 20 12
rect 26 -57 29 1
rect 34 -62 37 12
rect 42 -62 45 12
rect 50 -62 53 12
rect 58 -62 61 12
rect 66 -62 69 12
rect 74 -62 77 12
rect 82 -62 85 12
rect 90 -62 93 12
rect 98 -62 101 12
rect 106 -62 109 12
rect 277 9 280 22
rect 292 24 322 28
rect 292 19 296 24
rect 318 17 398 20
rect 314 9 317 16
rect 277 6 317 9
rect 326 6 396 10
rect 140 0 181 3
rect 196 0 215 3
rect 118 -4 132 -3
rect 118 -6 170 -4
rect 129 -7 170 -6
rect 178 -5 181 0
rect 281 -4 317 -1
rect 321 -4 408 -1
rect 178 -8 215 -5
rect 140 -16 181 -13
rect 249 -13 317 -10
rect 321 -12 408 -9
rect 196 -16 215 -13
rect 118 -20 132 -19
rect 118 -22 170 -20
rect 129 -23 170 -22
rect 178 -21 181 -16
rect 281 -20 317 -17
rect 321 -20 408 -17
rect 178 -24 215 -21
rect 140 -32 181 -29
rect 249 -29 317 -26
rect 321 -28 408 -25
rect 196 -32 215 -29
rect 118 -36 132 -35
rect 118 -38 170 -36
rect 129 -39 170 -38
rect 178 -37 181 -32
rect 281 -36 317 -33
rect 321 -36 408 -33
rect 178 -40 215 -37
rect 249 -45 317 -42
rect 321 -44 408 -41
rect 196 -48 215 -45
rect 118 -52 132 -51
rect 118 -54 170 -52
rect 129 -55 170 -54
rect 281 -52 317 -49
rect 321 -52 408 -49
rect 34 -65 38 -62
rect 42 -65 46 -62
rect 50 -65 54 -62
rect 58 -65 62 -62
rect 66 -65 70 -62
rect 74 -65 78 -62
rect 82 -65 86 -62
rect 90 -65 94 -62
rect 98 -65 102 -62
rect 106 -65 110 -62
rect 157 -64 292 -61
rect 35 -69 38 -65
rect 43 -69 46 -65
rect 51 -69 54 -65
rect 59 -69 62 -65
rect 67 -69 70 -65
rect 75 -69 78 -65
rect 83 -69 86 -65
rect 91 -69 94 -65
rect 99 -69 102 -65
rect 107 -69 110 -65
rect 120 -72 135 -69
rect 167 -72 177 -68
rect 181 -72 299 -68
rect 35 -114 38 -73
rect 43 -150 46 -73
rect 51 -114 54 -73
rect 59 -150 62 -73
rect 67 -114 70 -73
rect 75 -150 78 -73
rect 83 -114 86 -73
rect 91 -150 94 -73
rect 99 -114 102 -73
rect 107 -150 110 -73
rect 131 -80 208 -76
rect 212 -80 252 -76
rect 296 -86 323 -83
rect 120 -94 163 -90
rect 331 -95 334 -62
rect 347 -95 350 -62
rect 363 -95 366 -62
rect 379 -95 382 -62
rect 331 -98 343 -95
rect 347 -98 359 -95
rect 363 -98 375 -95
rect 379 -98 391 -95
rect 288 -138 323 -135
rect 43 -172 46 -154
rect 59 -172 62 -154
rect 75 -172 78 -154
rect 91 -172 94 -154
rect 107 -172 110 -154
rect 34 -175 46 -172
rect 50 -175 62 -172
rect 66 -175 78 -172
rect 82 -175 94 -172
rect 98 -175 110 -172
rect 5 -181 25 -177
rect 34 -189 37 -175
rect 50 -189 53 -175
rect 66 -189 69 -175
rect 82 -189 85 -175
rect 98 -189 101 -175
rect 131 -181 323 -177
rect 41 -197 44 -193
rect 57 -197 60 -193
rect 73 -197 76 -193
rect 89 -197 92 -193
rect 105 -197 108 -193
rect 12 -203 25 -200
rect 34 -200 44 -197
rect 50 -200 60 -197
rect 66 -200 76 -197
rect 82 -200 92 -197
rect 98 -200 108 -197
rect 5 -211 25 -207
rect 34 -221 37 -200
rect 12 -235 25 -232
rect 34 -273 37 -225
rect 42 -248 45 -218
rect 50 -221 53 -200
rect 42 -276 45 -252
rect 50 -273 53 -225
rect 58 -248 61 -218
rect 66 -221 69 -200
rect 58 -276 61 -252
rect 66 -273 69 -225
rect 74 -248 77 -218
rect 82 -221 85 -200
rect 74 -276 77 -252
rect 82 -273 85 -225
rect 90 -248 93 -218
rect 98 -221 101 -200
rect 120 -204 142 -201
rect 331 -205 334 -106
rect 340 -170 343 -98
rect 347 -205 350 -106
rect 356 -170 359 -98
rect 363 -205 366 -106
rect 372 -170 375 -98
rect 379 -205 382 -106
rect 388 -170 391 -98
rect 331 -208 342 -205
rect 347 -208 358 -205
rect 363 -208 374 -205
rect 379 -208 390 -205
rect 90 -276 93 -252
rect 98 -273 101 -225
rect 106 -248 109 -218
rect 120 -236 142 -233
rect 106 -276 109 -252
rect 296 -256 323 -253
rect 120 -265 135 -262
rect 331 -273 334 -236
rect 339 -273 342 -208
rect 347 -273 350 -236
rect 355 -273 358 -208
rect 363 -273 366 -236
rect 371 -273 374 -208
rect 379 -273 382 -236
rect 387 -273 390 -208
<< labels >>
rlabel metal2 42 -254 45 -254 1 RESET
rlabel metal2 58 -254 61 -254 1 load
rlabel metal2 74 -254 77 -254 1 iter
rlabel metal2 90 -254 93 -254 1 InSt0*
rlabel metal2 106 -254 109 -254 1 InSt1*
rlabel metal1 284 -272 287 -272 1 p1-
rlabel metal1 292 -272 295 -272 1 p1
rlabel metal1 143 -275 146 -275 1 p2-
rlabel metal1 135 -275 138 -275 1 p2
rlabel metal1 123 -275 131 -275 1 Vdd!
rlabel metal1 299 -272 307 -272 1 GND!
rlabel metal1 331 -230 334 -230 1 OutSt1*
rlabel metal2 339 -230 342 -230 1 OutSt0*
rlabel metal1 347 -230 350 -230 1 ready
rlabel metal2 355 -230 358 -230 1 sreg_en
rlabel metal1 363 -230 366 -230 1 sreg_latch
rlabel metal2 371 -230 374 -230 1 add_latch
rlabel metal1 379 -230 382 -230 1 in_latch
rlabel metal2 387 -230 390 -230 1 loop_latch
<< end >>
