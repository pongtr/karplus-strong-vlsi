magic
tech scmos
timestamp 1509371954
<< psubstratepdiff >>
rect 144 39 150 71
rect 159 39 165 71
<< metal1 >>
rect 97 356 213 357
rect 97 352 110 356
rect 114 352 117 356
rect 121 352 124 356
rect 128 352 131 356
rect 135 352 138 356
rect 142 352 145 356
rect 149 352 152 356
rect 156 352 159 356
rect 163 352 166 356
rect 170 352 173 356
rect 177 352 180 356
rect 184 352 187 356
rect 191 352 194 356
rect 198 352 213 356
rect 97 351 213 352
rect 97 348 110 351
rect 107 347 110 348
rect 114 347 117 351
rect 121 347 124 351
rect 128 347 131 351
rect 135 347 138 351
rect 142 347 145 351
rect 149 347 152 351
rect 156 347 159 351
rect 163 347 166 351
rect 170 347 173 351
rect 177 347 180 351
rect 184 347 187 351
rect 191 347 194 351
rect 198 348 213 351
rect 198 347 203 348
rect 107 346 203 347
rect 107 342 110 346
rect 114 342 117 346
rect 121 342 124 346
rect 128 342 131 346
rect 135 342 138 346
rect 142 342 145 346
rect 149 342 152 346
rect 156 342 159 346
rect 163 342 166 346
rect 170 342 173 346
rect 177 342 180 346
rect 184 342 187 346
rect 191 342 194 346
rect 198 342 203 346
rect 107 341 203 342
rect 107 337 110 341
rect 114 337 117 341
rect 121 337 124 341
rect 128 337 131 341
rect 135 337 138 341
rect 142 337 145 341
rect 149 337 152 341
rect 156 337 159 341
rect 163 337 166 341
rect 170 337 173 341
rect 177 337 180 341
rect 184 337 187 341
rect 191 337 194 341
rect 198 337 203 341
rect 107 336 203 337
rect 45 203 48 207
rect 52 203 53 207
rect 57 203 58 207
rect 62 203 63 207
rect 67 203 68 207
rect 72 203 73 207
rect 77 203 78 207
rect 82 203 83 207
rect 87 203 88 207
rect 92 203 93 207
rect 97 203 98 207
rect 102 203 105 207
rect 31 157 87 194
rect 19 155 87 157
rect 19 151 20 155
rect 24 151 25 155
rect 29 151 87 155
rect 19 150 87 151
rect 19 146 20 150
rect 24 146 25 150
rect 29 146 87 150
rect 19 145 87 146
rect 19 141 20 145
rect 24 141 25 145
rect 29 141 87 145
rect 19 140 87 141
rect 19 136 20 140
rect 24 136 25 140
rect 29 136 87 140
rect 19 135 87 136
rect 19 131 20 135
rect 24 131 25 135
rect 29 131 87 135
rect 19 130 87 131
rect 19 126 20 130
rect 24 126 25 130
rect 29 126 87 130
rect 19 125 87 126
rect 19 121 20 125
rect 24 121 25 125
rect 29 121 87 125
rect 19 120 87 121
rect 19 116 20 120
rect 24 116 25 120
rect 29 116 87 120
rect 19 115 87 116
rect 19 111 20 115
rect 24 111 25 115
rect 29 111 87 115
rect 19 110 87 111
rect 19 106 20 110
rect 24 106 25 110
rect 29 106 87 110
rect 19 105 87 106
rect 19 101 20 105
rect 24 101 25 105
rect 29 101 87 105
rect 19 100 87 101
rect 19 96 20 100
rect 24 96 25 100
rect 29 96 87 100
rect 19 95 87 96
rect 19 91 20 95
rect 24 91 25 95
rect 29 91 87 95
rect 19 89 87 91
rect 129 70 181 336
rect 205 203 208 207
rect 212 203 213 207
rect 217 203 218 207
rect 222 203 223 207
rect 227 203 228 207
rect 232 203 233 207
rect 237 203 238 207
rect 242 203 243 207
rect 247 203 248 207
rect 252 203 253 207
rect 257 203 258 207
rect 262 203 265 207
rect 129 66 155 70
rect 159 66 160 70
rect 164 66 181 70
rect 225 77 281 194
rect 229 73 230 77
rect 234 73 235 77
rect 239 73 240 77
rect 244 73 245 77
rect 249 73 250 77
rect 254 73 255 77
rect 259 73 260 77
rect 264 73 265 77
rect 269 73 270 77
rect 274 73 275 77
rect 279 73 281 77
rect 225 72 281 73
rect 229 68 230 72
rect 234 68 235 72
rect 239 68 240 72
rect 244 68 245 72
rect 249 68 250 72
rect 254 68 255 72
rect 259 68 260 72
rect 264 68 265 72
rect 269 68 270 72
rect 274 68 275 72
rect 279 68 281 72
rect 225 67 281 68
rect 129 65 181 66
rect 129 61 155 65
rect 159 61 160 65
rect 164 61 181 65
rect 129 60 181 61
rect 129 56 155 60
rect 159 56 160 60
rect 164 56 181 60
rect 129 55 181 56
rect 129 51 155 55
rect 159 51 160 55
rect 164 51 181 55
rect 129 50 181 51
rect 129 46 155 50
rect 159 46 160 50
rect 164 46 181 50
rect 129 45 181 46
rect 129 41 155 45
rect 159 41 160 45
rect 164 41 181 45
rect 129 40 181 41
rect 129 36 155 40
rect 159 36 160 40
rect 164 36 181 40
rect 129 35 181 36
rect 129 31 155 35
rect 159 31 160 35
rect 164 31 181 35
rect 129 30 181 31
rect 129 26 155 30
rect 159 26 160 30
rect 164 26 181 30
rect 129 25 181 26
rect 129 21 155 25
rect 159 21 160 25
rect 164 21 181 25
rect 129 20 181 21
rect 129 16 155 20
rect 159 16 160 20
rect 164 16 181 20
rect 129 -35 181 16
<< m2contact >>
rect 110 352 114 356
rect 117 352 121 356
rect 124 352 128 356
rect 131 352 135 356
rect 138 352 142 356
rect 145 352 149 356
rect 152 352 156 356
rect 159 352 163 356
rect 166 352 170 356
rect 173 352 177 356
rect 180 352 184 356
rect 187 352 191 356
rect 194 352 198 356
rect 110 347 114 351
rect 117 347 121 351
rect 124 347 128 351
rect 131 347 135 351
rect 138 347 142 351
rect 145 347 149 351
rect 152 347 156 351
rect 159 347 163 351
rect 166 347 170 351
rect 173 347 177 351
rect 180 347 184 351
rect 187 347 191 351
rect 194 347 198 351
rect 110 342 114 346
rect 117 342 121 346
rect 124 342 128 346
rect 131 342 135 346
rect 138 342 142 346
rect 145 342 149 346
rect 152 342 156 346
rect 159 342 163 346
rect 166 342 170 346
rect 173 342 177 346
rect 180 342 184 346
rect 187 342 191 346
rect 194 342 198 346
rect 110 337 114 341
rect 117 337 121 341
rect 124 337 128 341
rect 131 337 135 341
rect 138 337 142 341
rect 145 337 149 341
rect 152 337 156 341
rect 159 337 163 341
rect 166 337 170 341
rect 173 337 177 341
rect 180 337 184 341
rect 187 337 191 341
rect 194 337 198 341
rect 41 203 45 207
rect 48 203 52 207
rect 53 203 57 207
rect 58 203 62 207
rect 63 203 67 207
rect 68 203 72 207
rect 73 203 77 207
rect 78 203 82 207
rect 83 203 87 207
rect 88 203 92 207
rect 93 203 97 207
rect 98 203 102 207
rect 105 203 109 207
rect 20 151 24 155
rect 25 151 29 155
rect 20 146 24 150
rect 25 146 29 150
rect 20 141 24 145
rect 25 141 29 145
rect 20 136 24 140
rect 25 136 29 140
rect 20 131 24 135
rect 25 131 29 135
rect 20 126 24 130
rect 25 126 29 130
rect 20 121 24 125
rect 25 121 29 125
rect 20 116 24 120
rect 25 116 29 120
rect 20 111 24 115
rect 25 111 29 115
rect 20 106 24 110
rect 25 106 29 110
rect 20 101 24 105
rect 25 101 29 105
rect 20 96 24 100
rect 25 96 29 100
rect 20 91 24 95
rect 25 91 29 95
rect 201 203 205 207
rect 208 203 212 207
rect 213 203 217 207
rect 218 203 222 207
rect 223 203 227 207
rect 228 203 232 207
rect 233 203 237 207
rect 238 203 242 207
rect 243 203 247 207
rect 248 203 252 207
rect 253 203 257 207
rect 258 203 262 207
rect 265 203 269 207
rect 155 66 159 70
rect 160 66 164 70
rect 225 73 229 77
rect 230 73 234 77
rect 235 73 239 77
rect 240 73 244 77
rect 245 73 249 77
rect 250 73 254 77
rect 255 73 259 77
rect 260 73 264 77
rect 265 73 269 77
rect 270 73 274 77
rect 275 73 279 77
rect 225 68 229 72
rect 230 68 234 72
rect 235 68 239 72
rect 240 68 244 72
rect 245 68 249 72
rect 250 68 254 72
rect 255 68 259 72
rect 260 68 264 72
rect 265 68 269 72
rect 270 68 274 72
rect 275 68 279 72
rect 155 61 159 65
rect 160 61 164 65
rect 155 56 159 60
rect 160 56 164 60
rect 155 51 159 55
rect 160 51 164 55
rect 155 46 159 50
rect 160 46 164 50
rect 155 41 159 45
rect 160 41 164 45
rect 155 36 159 40
rect 160 36 164 40
rect 155 31 159 35
rect 160 31 164 35
rect 155 26 159 30
rect 160 26 164 30
rect 155 21 159 25
rect 160 21 164 25
rect 155 16 159 20
rect 160 16 164 20
<< metal2 >>
rect 97 356 213 357
rect 97 352 110 356
rect 114 352 117 356
rect 121 352 124 356
rect 128 352 131 356
rect 135 352 138 356
rect 142 352 145 356
rect 149 352 152 356
rect 156 352 159 356
rect 163 352 166 356
rect 170 352 173 356
rect 177 352 180 356
rect 184 352 187 356
rect 191 352 194 356
rect 198 352 213 356
rect 97 351 213 352
rect 97 348 110 351
rect 107 347 110 348
rect 114 347 117 351
rect 121 347 124 351
rect 128 347 131 351
rect 135 347 138 351
rect 142 347 145 351
rect 149 347 152 351
rect 156 347 159 351
rect 163 347 166 351
rect 170 347 173 351
rect 177 347 180 351
rect 184 347 187 351
rect 191 347 194 351
rect 198 348 213 351
rect 198 347 203 348
rect 107 346 203 347
rect 107 342 110 346
rect 114 342 117 346
rect 121 342 124 346
rect 128 342 131 346
rect 135 342 138 346
rect 142 342 145 346
rect 149 342 152 346
rect 156 342 159 346
rect 163 342 166 346
rect 170 342 173 346
rect 177 342 180 346
rect 184 342 187 346
rect 191 342 194 346
rect 198 342 203 346
rect 107 341 203 342
rect 107 337 110 341
rect 114 337 117 341
rect 121 337 124 341
rect 128 337 131 341
rect 135 337 138 341
rect 142 337 145 341
rect 149 337 152 341
rect 156 337 159 341
rect 163 337 166 341
rect 170 337 173 341
rect 177 337 180 341
rect 184 337 187 341
rect 191 337 194 341
rect 198 337 203 341
rect 107 308 203 337
rect 97 219 213 308
rect 45 203 48 207
rect 52 203 53 207
rect 57 203 58 207
rect 62 203 63 207
rect 67 203 68 207
rect 72 203 73 207
rect 77 203 78 207
rect 82 203 83 207
rect 87 203 88 207
rect 92 203 93 207
rect 97 203 98 207
rect 102 203 105 207
rect 8 155 29 157
rect 8 151 10 155
rect 14 151 15 155
rect 19 151 20 155
rect 24 151 25 155
rect 8 150 29 151
rect 8 146 10 150
rect 14 146 15 150
rect 19 146 20 150
rect 24 146 25 150
rect 8 145 29 146
rect 8 141 10 145
rect 14 141 15 145
rect 19 141 20 145
rect 24 141 25 145
rect 8 140 29 141
rect 8 136 10 140
rect 14 136 15 140
rect 19 136 20 140
rect 24 136 25 140
rect 8 135 29 136
rect 8 131 10 135
rect 14 131 15 135
rect 19 131 20 135
rect 24 131 25 135
rect 8 130 29 131
rect 8 126 10 130
rect 14 126 15 130
rect 19 126 20 130
rect 24 126 25 130
rect 8 125 29 126
rect 8 121 10 125
rect 14 121 15 125
rect 19 121 20 125
rect 24 121 25 125
rect 8 120 29 121
rect 8 116 10 120
rect 14 116 15 120
rect 19 116 20 120
rect 24 116 25 120
rect 8 115 29 116
rect 8 111 10 115
rect 14 111 15 115
rect 19 111 20 115
rect 24 111 25 115
rect 8 110 29 111
rect 8 106 10 110
rect 14 106 15 110
rect 19 106 20 110
rect 24 106 25 110
rect 8 105 29 106
rect 8 101 10 105
rect 14 101 15 105
rect 19 101 20 105
rect 24 101 25 105
rect 8 100 29 101
rect 8 96 10 100
rect 14 96 15 100
rect 19 96 20 100
rect 24 96 25 100
rect 8 95 29 96
rect 8 91 10 95
rect 14 91 15 95
rect 19 91 20 95
rect 24 91 25 95
rect 8 89 29 91
rect 41 67 109 203
rect 205 203 208 207
rect 212 203 213 207
rect 217 203 218 207
rect 222 203 223 207
rect 227 203 228 207
rect 232 203 233 207
rect 237 203 238 207
rect 242 203 243 207
rect 247 203 248 207
rect 252 203 253 207
rect 257 203 258 207
rect 262 203 265 207
rect 201 124 269 203
rect 201 120 203 124
rect 207 120 208 124
rect 212 120 213 124
rect 217 120 218 124
rect 222 120 223 124
rect 227 120 228 124
rect 232 120 233 124
rect 237 120 238 124
rect 242 120 243 124
rect 247 120 248 124
rect 252 120 253 124
rect 257 120 258 124
rect 262 120 263 124
rect 267 120 269 124
rect 201 119 269 120
rect 201 115 203 119
rect 207 115 208 119
rect 212 115 213 119
rect 217 115 218 119
rect 222 115 223 119
rect 227 115 228 119
rect 232 115 233 119
rect 237 115 238 119
rect 242 115 243 119
rect 247 115 248 119
rect 252 115 253 119
rect 257 115 258 119
rect 262 115 263 119
rect 267 115 269 119
rect 201 112 269 115
rect 229 73 230 77
rect 234 73 235 77
rect 239 73 240 77
rect 244 73 245 77
rect 249 73 250 77
rect 254 73 255 77
rect 259 73 260 77
rect 264 73 265 77
rect 269 73 270 77
rect 274 73 275 77
rect 279 73 281 77
rect 225 72 281 73
rect 41 63 43 67
rect 47 63 48 67
rect 52 63 53 67
rect 57 63 58 67
rect 62 63 63 67
rect 67 63 68 67
rect 72 63 73 67
rect 77 63 78 67
rect 82 63 83 67
rect 87 63 88 67
rect 92 63 93 67
rect 97 63 98 67
rect 102 63 103 67
rect 107 63 109 67
rect 41 62 109 63
rect 41 58 43 62
rect 47 58 48 62
rect 52 58 53 62
rect 57 58 58 62
rect 62 58 63 62
rect 67 58 68 62
rect 72 58 73 62
rect 77 58 78 62
rect 82 58 83 62
rect 87 58 88 62
rect 92 58 93 62
rect 97 58 98 62
rect 102 58 103 62
rect 107 58 109 62
rect 41 55 109 58
rect 144 66 145 70
rect 149 66 150 70
rect 154 66 155 70
rect 159 66 160 70
rect 144 65 164 66
rect 144 61 145 65
rect 149 61 150 65
rect 154 61 155 65
rect 159 61 160 65
rect 144 60 164 61
rect 144 56 145 60
rect 149 56 150 60
rect 154 56 155 60
rect 159 56 160 60
rect 229 68 230 72
rect 234 68 235 72
rect 239 68 240 72
rect 244 68 245 72
rect 249 68 250 72
rect 254 68 255 72
rect 259 68 260 72
rect 264 68 265 72
rect 269 68 270 72
rect 274 68 275 72
rect 279 68 281 72
rect 225 67 281 68
rect 229 63 230 67
rect 234 63 235 67
rect 239 63 240 67
rect 244 63 245 67
rect 249 63 250 67
rect 254 63 255 67
rect 259 63 260 67
rect 264 63 265 67
rect 269 63 270 67
rect 274 63 275 67
rect 279 63 281 67
rect 225 62 281 63
rect 229 58 230 62
rect 234 58 235 62
rect 239 58 240 62
rect 244 58 245 62
rect 249 58 250 62
rect 254 58 255 62
rect 259 58 260 62
rect 264 58 265 62
rect 269 58 270 62
rect 274 58 275 62
rect 279 58 281 62
rect 225 56 281 58
rect 144 55 164 56
rect 144 51 145 55
rect 149 51 150 55
rect 154 51 155 55
rect 159 51 160 55
rect 144 50 164 51
rect 144 46 145 50
rect 149 46 150 50
rect 154 46 155 50
rect 159 46 160 50
rect 144 45 164 46
rect 144 41 145 45
rect 149 41 150 45
rect 154 41 155 45
rect 159 41 160 45
rect 144 40 164 41
rect 144 36 145 40
rect 149 36 150 40
rect 154 36 155 40
rect 159 36 160 40
rect 144 35 164 36
rect 144 31 145 35
rect 149 31 150 35
rect 154 31 155 35
rect 159 31 160 35
rect 144 30 164 31
rect 144 26 145 30
rect 149 26 150 30
rect 154 26 155 30
rect 159 26 160 30
rect 144 25 164 26
rect 144 21 145 25
rect 149 21 150 25
rect 154 21 155 25
rect 159 21 160 25
rect 144 20 164 21
rect 144 16 145 20
rect 149 16 150 20
rect 154 16 155 20
rect 159 16 160 20
rect 144 14 164 16
<< m3contact >>
rect 10 151 14 155
rect 15 151 19 155
rect 10 146 14 150
rect 15 146 19 150
rect 10 141 14 145
rect 15 141 19 145
rect 10 136 14 140
rect 15 136 19 140
rect 10 131 14 135
rect 15 131 19 135
rect 10 126 14 130
rect 15 126 19 130
rect 10 121 14 125
rect 15 121 19 125
rect 10 116 14 120
rect 15 116 19 120
rect 10 111 14 115
rect 15 111 19 115
rect 10 106 14 110
rect 15 106 19 110
rect 10 101 14 105
rect 15 101 19 105
rect 10 96 14 100
rect 15 96 19 100
rect 10 91 14 95
rect 15 91 19 95
rect 203 120 207 124
rect 208 120 212 124
rect 213 120 217 124
rect 218 120 222 124
rect 223 120 227 124
rect 228 120 232 124
rect 233 120 237 124
rect 238 120 242 124
rect 243 120 247 124
rect 248 120 252 124
rect 253 120 257 124
rect 258 120 262 124
rect 263 120 267 124
rect 203 115 207 119
rect 208 115 212 119
rect 213 115 217 119
rect 218 115 222 119
rect 223 115 227 119
rect 228 115 232 119
rect 233 115 237 119
rect 238 115 242 119
rect 243 115 247 119
rect 248 115 252 119
rect 253 115 257 119
rect 258 115 262 119
rect 263 115 267 119
rect 43 63 47 67
rect 48 63 52 67
rect 53 63 57 67
rect 58 63 62 67
rect 63 63 67 67
rect 68 63 72 67
rect 73 63 77 67
rect 78 63 82 67
rect 83 63 87 67
rect 88 63 92 67
rect 93 63 97 67
rect 98 63 102 67
rect 103 63 107 67
rect 43 58 47 62
rect 48 58 52 62
rect 53 58 57 62
rect 58 58 62 62
rect 63 58 67 62
rect 68 58 72 62
rect 73 58 77 62
rect 78 58 82 62
rect 83 58 87 62
rect 88 58 92 62
rect 93 58 97 62
rect 98 58 102 62
rect 103 58 107 62
rect 145 66 149 70
rect 150 66 154 70
rect 145 61 149 65
rect 150 61 154 65
rect 145 56 149 60
rect 150 56 154 60
rect 225 63 229 67
rect 230 63 234 67
rect 235 63 239 67
rect 240 63 244 67
rect 245 63 249 67
rect 250 63 254 67
rect 255 63 259 67
rect 260 63 264 67
rect 265 63 269 67
rect 270 63 274 67
rect 275 63 279 67
rect 225 58 229 62
rect 230 58 234 62
rect 235 58 239 62
rect 240 58 244 62
rect 245 58 249 62
rect 250 58 254 62
rect 255 58 259 62
rect 260 58 264 62
rect 265 58 269 62
rect 270 58 274 62
rect 275 58 279 62
rect 145 51 149 55
rect 150 51 154 55
rect 145 46 149 50
rect 150 46 154 50
rect 145 41 149 45
rect 150 41 154 45
rect 145 36 149 40
rect 150 36 154 40
rect 145 31 149 35
rect 150 31 154 35
rect 145 26 149 30
rect 150 26 154 30
rect 145 21 149 25
rect 150 21 154 25
rect 145 16 149 20
rect 150 16 154 20
<< metal3 >>
rect 8 155 20 157
rect 8 151 10 155
rect 14 151 15 155
rect 19 151 20 155
rect 8 150 20 151
rect 8 146 10 150
rect 14 146 15 150
rect 19 146 20 150
rect 8 145 20 146
rect 8 141 10 145
rect 14 141 15 145
rect 19 141 20 145
rect 8 140 20 141
rect 8 136 10 140
rect 14 136 15 140
rect 19 136 20 140
rect 8 135 20 136
rect 8 131 10 135
rect 14 131 15 135
rect 19 131 20 135
rect 8 130 20 131
rect 8 126 10 130
rect 14 126 15 130
rect 19 126 20 130
rect 8 125 20 126
rect 8 121 10 125
rect 14 121 15 125
rect 19 121 20 125
rect 8 120 20 121
rect 8 116 10 120
rect 14 116 15 120
rect 19 116 20 120
rect 8 115 20 116
rect 8 111 10 115
rect 14 111 15 115
rect 19 111 20 115
rect 201 124 269 125
rect 201 120 203 124
rect 207 120 208 124
rect 212 120 213 124
rect 217 120 218 124
rect 222 120 223 124
rect 227 120 228 124
rect 232 120 233 124
rect 237 120 238 124
rect 242 120 243 124
rect 247 120 248 124
rect 252 120 253 124
rect 257 120 258 124
rect 262 120 263 124
rect 267 120 269 124
rect 201 119 269 120
rect 201 115 203 119
rect 207 115 208 119
rect 212 115 213 119
rect 217 115 218 119
rect 222 115 223 119
rect 227 115 228 119
rect 232 115 233 119
rect 237 115 238 119
rect 242 115 243 119
rect 247 115 248 119
rect 252 115 253 119
rect 257 115 258 119
rect 262 115 263 119
rect 267 115 269 119
rect 201 112 269 115
rect 8 110 20 111
rect 8 106 10 110
rect 14 106 15 110
rect 19 106 20 110
rect 8 105 20 106
rect 8 101 10 105
rect 14 101 15 105
rect 19 101 20 105
rect 8 100 20 101
rect 8 96 10 100
rect 14 96 15 100
rect 19 96 20 100
rect 8 95 20 96
rect 8 91 10 95
rect 14 91 15 95
rect 19 91 20 95
rect 8 88 20 91
rect 144 70 165 71
rect 41 67 109 68
rect 41 63 43 67
rect 47 63 48 67
rect 52 63 53 67
rect 57 63 58 67
rect 62 63 63 67
rect 67 63 68 67
rect 72 63 73 67
rect 77 63 78 67
rect 82 63 83 67
rect 87 63 88 67
rect 92 63 93 67
rect 97 63 98 67
rect 102 63 103 67
rect 107 63 109 67
rect 41 62 109 63
rect 41 58 43 62
rect 47 58 48 62
rect 52 58 53 62
rect 57 58 58 62
rect 62 58 63 62
rect 67 58 68 62
rect 72 58 73 62
rect 77 58 78 62
rect 82 58 83 62
rect 87 58 88 62
rect 92 58 93 62
rect 97 58 98 62
rect 102 58 103 62
rect 107 58 109 62
rect 41 55 109 58
rect 144 66 145 70
rect 149 66 150 70
rect 154 66 165 70
rect 144 65 165 66
rect 144 61 145 65
rect 149 61 150 65
rect 154 61 165 65
rect 144 60 165 61
rect 144 56 145 60
rect 149 56 150 60
rect 154 56 165 60
rect 224 67 281 69
rect 224 63 225 67
rect 229 63 230 67
rect 234 63 235 67
rect 239 63 240 67
rect 244 63 245 67
rect 249 63 250 67
rect 254 63 255 67
rect 259 63 260 67
rect 264 63 265 67
rect 269 63 270 67
rect 274 63 275 67
rect 279 63 281 67
rect 224 62 281 63
rect 224 58 225 62
rect 229 58 230 62
rect 234 58 235 62
rect 239 58 240 62
rect 244 58 245 62
rect 249 58 250 62
rect 254 58 255 62
rect 259 58 260 62
rect 264 58 265 62
rect 269 58 270 62
rect 274 58 275 62
rect 279 58 281 62
rect 224 56 281 58
rect 144 55 165 56
rect 144 51 145 55
rect 149 51 150 55
rect 154 51 165 55
rect 144 50 165 51
rect 144 46 145 50
rect 149 46 150 50
rect 154 46 165 50
rect 144 45 165 46
rect 144 41 145 45
rect 149 41 150 45
rect 154 41 165 45
rect 144 40 165 41
rect 144 36 145 40
rect 149 36 150 40
rect 154 36 165 40
rect 144 35 165 36
rect 144 31 145 35
rect 149 31 150 35
rect 154 31 165 35
rect 144 30 165 31
rect 144 26 145 30
rect 149 26 150 30
rect 154 26 165 30
rect 144 25 165 26
rect 144 21 145 25
rect 149 21 150 25
rect 154 21 165 25
rect 144 20 165 21
rect 144 16 145 20
rect 149 16 150 20
rect 154 16 165 20
rect 144 14 165 16
use barepad  b
timestamp 1006127261
transform 1 0 9 0 1 -366
box 16 702 276 1014
use ndiode  nd
timestamp 1037203521
transform 1 0 41 0 1 206
box -14 -13 82 128
use pdiode  pd
timestamp 1037203492
transform 1 0 180 0 1 202
box 7 -9 103 132
use barering  br
timestamp 1006127261
transform 1 0 -2 0 1 -12
box 2 -23 311 176
<< labels >>
rlabel metal3 15 94 15 94 1 Vdd!
rlabel metal1 153 210 153 210 1 GND!
<< end >>
