magic
tech scmos
timestamp 1512683628
<< checkpaint >>
rect -1 -286 413 34
<< polysilicon >>
rect 324 21 331 23
rect 335 21 339 23
rect 343 21 347 23
rect 351 21 355 23
rect 359 21 363 23
rect 367 21 371 23
rect 375 21 379 23
rect 383 21 387 23
rect 391 21 398 23
rect 10 -2 12 3
rect 10 -10 12 -6
rect 10 -18 12 -14
rect 10 -26 12 -22
rect 10 -34 12 -30
rect 10 -42 12 -38
rect 10 -50 12 -46
rect 10 -58 12 -54
rect 10 -67 12 -62
rect 34 -72 36 8
rect 42 -50 44 8
rect 42 -58 44 -54
rect 50 -58 52 8
rect 42 -72 44 -62
rect 50 -72 52 -62
rect 58 -72 60 8
rect 66 -50 68 8
rect 66 -72 68 -54
rect 74 -72 76 8
rect 82 -26 84 8
rect 90 -2 92 8
rect 90 -10 92 -6
rect 98 -10 100 8
rect 106 -2 108 8
rect 127 5 129 7
rect 133 5 145 7
rect 149 5 152 7
rect 156 5 185 7
rect 189 5 201 7
rect 205 5 207 7
rect 119 -3 129 -1
rect 133 -3 156 -1
rect 160 -3 162 -1
rect 223 0 254 2
rect 274 0 286 2
rect 296 0 298 2
rect 174 -3 177 -1
rect 181 -3 201 -1
rect 205 -3 207 -1
rect 82 -34 84 -30
rect 82 -42 84 -38
rect 82 -72 84 -46
rect 90 -72 92 -14
rect 98 -18 100 -14
rect 98 -72 100 -22
rect 106 -26 108 -6
rect 119 -12 121 -3
rect 127 -11 129 -9
rect 133 -11 145 -9
rect 149 -11 152 -9
rect 326 -3 347 -1
rect 351 -3 403 -1
rect 223 -8 224 -6
rect 244 -8 306 -6
rect 316 -8 318 -6
rect 156 -11 185 -9
rect 189 -11 201 -9
rect 205 -11 207 -9
rect 119 -19 129 -17
rect 133 -19 156 -17
rect 160 -19 162 -17
rect 326 -11 355 -9
rect 359 -11 363 -9
rect 367 -11 403 -9
rect 223 -16 254 -14
rect 274 -16 286 -14
rect 296 -16 298 -14
rect 174 -19 177 -17
rect 181 -19 201 -17
rect 205 -19 207 -17
rect 119 -28 121 -19
rect 127 -27 129 -25
rect 133 -27 145 -25
rect 149 -27 152 -25
rect 106 -72 108 -30
rect 326 -19 379 -17
rect 383 -19 403 -17
rect 223 -24 224 -22
rect 244 -24 306 -22
rect 316 -24 318 -22
rect 156 -27 185 -25
rect 189 -27 201 -25
rect 205 -27 207 -25
rect 119 -35 129 -33
rect 133 -35 156 -33
rect 160 -35 162 -33
rect 326 -27 387 -25
rect 391 -27 403 -25
rect 223 -32 254 -30
rect 274 -32 286 -30
rect 296 -32 298 -30
rect 174 -35 177 -33
rect 181 -35 201 -33
rect 205 -35 207 -33
rect 119 -44 121 -35
rect 127 -43 129 -41
rect 133 -43 145 -41
rect 149 -43 152 -41
rect 326 -35 355 -33
rect 359 -35 403 -33
rect 223 -40 224 -38
rect 244 -40 306 -38
rect 316 -40 318 -38
rect 156 -43 185 -41
rect 189 -43 201 -41
rect 205 -43 207 -41
rect 119 -51 129 -49
rect 133 -51 156 -49
rect 160 -51 162 -49
rect 326 -43 371 -41
rect 375 -43 403 -41
rect 223 -48 254 -46
rect 274 -48 286 -46
rect 296 -48 298 -46
rect 174 -51 177 -49
rect 181 -51 201 -49
rect 205 -51 207 -49
rect 119 -60 121 -51
rect 326 -51 339 -49
rect 343 -51 403 -49
rect 223 -56 224 -54
rect 244 -56 306 -54
rect 316 -56 318 -54
rect 326 -59 331 -57
rect 335 -59 403 -57
rect 343 -70 346 -68
rect 359 -70 362 -68
rect 375 -70 378 -68
rect 391 -70 394 -68
rect 344 -80 346 -70
rect 40 -82 42 -80
rect 56 -82 58 -80
rect 72 -82 74 -80
rect 88 -82 90 -80
rect 104 -82 106 -80
rect 32 -105 34 -103
rect 32 -130 34 -118
rect 32 -192 34 -155
rect 40 -165 42 -95
rect 48 -105 50 -103
rect 48 -130 50 -118
rect 40 -192 42 -191
rect 48 -192 50 -155
rect 56 -165 58 -95
rect 64 -105 66 -103
rect 64 -130 66 -118
rect 56 -192 58 -191
rect 64 -192 66 -155
rect 72 -165 74 -95
rect 80 -105 82 -103
rect 80 -130 82 -118
rect 72 -192 74 -191
rect 80 -192 82 -155
rect 88 -165 90 -95
rect 360 -80 362 -70
rect 336 -95 338 -94
rect 96 -105 98 -103
rect 96 -130 98 -118
rect 88 -192 90 -191
rect 96 -192 98 -155
rect 104 -165 106 -95
rect 336 -109 338 -105
rect 336 -117 338 -115
rect 336 -142 338 -141
rect 344 -144 346 -92
rect 376 -80 378 -70
rect 352 -95 354 -94
rect 352 -109 354 -105
rect 352 -117 354 -115
rect 352 -142 354 -141
rect 104 -192 106 -191
rect 39 -208 41 -207
rect 36 -209 41 -208
rect 45 -209 47 -207
rect 55 -208 57 -207
rect 52 -209 57 -208
rect 61 -209 63 -207
rect 71 -208 73 -207
rect 68 -209 73 -208
rect 77 -209 79 -207
rect 87 -208 89 -207
rect 84 -209 89 -208
rect 93 -209 95 -207
rect 103 -208 105 -207
rect 100 -209 105 -208
rect 109 -209 111 -207
rect 38 -214 41 -212
rect 45 -214 47 -212
rect 54 -214 57 -212
rect 61 -214 63 -212
rect 70 -214 73 -212
rect 77 -214 79 -212
rect 86 -214 89 -212
rect 93 -214 95 -212
rect 102 -214 105 -212
rect 109 -214 111 -212
rect 336 -213 338 -146
rect 360 -144 362 -92
rect 392 -80 394 -70
rect 368 -95 370 -94
rect 368 -109 370 -105
rect 368 -117 370 -115
rect 368 -142 370 -141
rect 344 -170 346 -168
rect 344 -185 346 -182
rect 38 -222 40 -214
rect 54 -222 56 -214
rect 70 -222 72 -214
rect 86 -222 88 -214
rect 102 -222 104 -214
rect 39 -240 41 -239
rect 36 -241 41 -240
rect 45 -241 47 -239
rect 55 -240 57 -239
rect 52 -241 57 -240
rect 61 -241 63 -239
rect 71 -240 73 -239
rect 68 -241 73 -240
rect 77 -241 79 -239
rect 87 -240 89 -239
rect 84 -241 89 -240
rect 93 -241 95 -239
rect 336 -239 338 -235
rect 103 -240 105 -239
rect 100 -241 105 -240
rect 109 -241 111 -239
rect 38 -246 41 -244
rect 45 -246 47 -244
rect 54 -246 57 -244
rect 61 -246 63 -244
rect 70 -246 73 -244
rect 77 -246 79 -244
rect 86 -246 89 -244
rect 93 -246 95 -244
rect 102 -246 105 -244
rect 109 -246 111 -244
rect 38 -256 40 -246
rect 54 -256 56 -246
rect 70 -256 72 -246
rect 86 -256 88 -246
rect 102 -256 104 -246
rect 336 -247 338 -245
rect 336 -260 338 -259
rect 38 -268 40 -260
rect 54 -268 56 -260
rect 70 -268 72 -260
rect 86 -268 88 -260
rect 102 -268 104 -260
rect 344 -262 346 -209
rect 352 -213 354 -146
rect 376 -144 378 -92
rect 384 -95 386 -94
rect 384 -109 386 -105
rect 384 -117 386 -115
rect 384 -142 386 -141
rect 360 -170 362 -168
rect 360 -185 362 -182
rect 352 -239 354 -235
rect 352 -247 354 -245
rect 352 -260 354 -259
rect 38 -270 41 -268
rect 45 -270 47 -268
rect 54 -270 57 -268
rect 61 -270 63 -268
rect 70 -270 73 -268
rect 77 -270 79 -268
rect 86 -270 89 -268
rect 93 -270 95 -268
rect 102 -270 105 -268
rect 109 -270 111 -268
rect 37 -274 41 -273
rect 39 -275 41 -274
rect 45 -275 47 -273
rect 53 -274 57 -273
rect 55 -275 57 -274
rect 61 -275 63 -273
rect 69 -274 73 -273
rect 71 -275 73 -274
rect 77 -275 79 -273
rect 85 -274 89 -273
rect 87 -275 89 -274
rect 93 -275 95 -273
rect 101 -274 105 -273
rect 103 -275 105 -274
rect 109 -275 111 -273
rect 360 -262 362 -209
rect 368 -213 370 -146
rect 392 -144 394 -92
rect 376 -170 378 -168
rect 376 -185 378 -182
rect 368 -239 370 -235
rect 368 -247 370 -245
rect 368 -260 370 -259
rect 344 -276 346 -274
rect 376 -262 378 -209
rect 384 -213 386 -146
rect 392 -170 394 -168
rect 392 -185 394 -182
rect 384 -239 386 -235
rect 384 -247 386 -245
rect 384 -260 386 -259
rect 360 -276 362 -274
rect 392 -262 394 -209
rect 376 -276 378 -274
rect 392 -276 394 -274
<< ndiffusion >>
rect 37 -50 41 1
rect 37 -54 42 -50
rect 44 -54 45 -50
rect 37 -58 41 -54
rect 53 -58 57 1
rect 37 -62 42 -58
rect 44 -62 45 -58
rect 49 -62 50 -58
rect 52 -62 57 -58
rect 37 -65 41 -62
rect 53 -65 57 -62
rect 69 -50 73 1
rect 65 -54 66 -50
rect 68 -54 73 -50
rect 69 -65 73 -54
rect 85 -2 89 1
rect 85 -6 90 -2
rect 92 -6 93 -2
rect 85 -10 89 -6
rect 101 -2 105 1
rect 145 7 149 8
rect 145 3 149 5
rect 185 7 189 8
rect 185 3 189 5
rect 145 0 160 3
rect 156 -1 160 0
rect 101 -6 106 -2
rect 108 -6 109 -2
rect 177 0 189 3
rect 177 -1 181 0
rect 286 2 296 3
rect 101 -10 105 -6
rect 85 -14 90 -10
rect 92 -14 93 -10
rect 97 -14 98 -10
rect 100 -14 105 -10
rect 85 -26 89 -14
rect 81 -30 82 -26
rect 84 -30 89 -26
rect 85 -34 89 -30
rect 81 -38 82 -34
rect 84 -38 89 -34
rect 85 -42 89 -38
rect 81 -46 82 -42
rect 84 -46 89 -42
rect 85 -65 89 -46
rect 101 -18 105 -14
rect 97 -22 98 -18
rect 100 -22 105 -18
rect 101 -26 105 -22
rect 156 -4 160 -3
rect 177 -4 181 -3
rect 156 -7 159 -4
rect 145 -9 149 -8
rect 145 -13 149 -11
rect 185 -9 189 -8
rect 286 -1 296 0
rect 347 -1 351 0
rect 298 -5 299 -1
rect 303 -5 304 -1
rect 314 -5 316 -1
rect 347 -4 351 -3
rect 306 -6 316 -5
rect 327 -8 396 -4
rect 306 -9 316 -8
rect 355 -9 359 -8
rect 363 -9 367 -8
rect 185 -13 189 -11
rect 145 -16 160 -13
rect 156 -17 160 -16
rect 177 -16 189 -13
rect 177 -17 181 -16
rect 355 -12 359 -11
rect 286 -14 296 -13
rect 363 -12 367 -11
rect 101 -30 106 -26
rect 108 -30 109 -26
rect 156 -20 160 -19
rect 177 -20 181 -19
rect 156 -23 159 -20
rect 145 -25 149 -24
rect 101 -65 105 -30
rect 145 -29 149 -27
rect 185 -25 189 -24
rect 286 -17 296 -16
rect 379 -17 383 -16
rect 298 -21 299 -17
rect 303 -21 304 -17
rect 314 -21 316 -17
rect 379 -20 383 -19
rect 306 -22 316 -21
rect 327 -24 396 -20
rect 306 -25 316 -24
rect 387 -25 391 -24
rect 185 -29 189 -27
rect 145 -32 160 -29
rect 156 -33 160 -32
rect 177 -32 189 -29
rect 177 -33 181 -32
rect 387 -28 391 -27
rect 286 -30 296 -29
rect 156 -36 160 -35
rect 177 -36 181 -35
rect 156 -39 159 -36
rect 145 -41 149 -40
rect 145 -45 149 -43
rect 185 -41 189 -40
rect 286 -33 296 -32
rect 355 -33 359 -32
rect 298 -37 299 -33
rect 303 -37 304 -33
rect 314 -37 316 -33
rect 355 -36 359 -35
rect 306 -38 316 -37
rect 327 -40 396 -36
rect 306 -41 316 -40
rect 371 -41 375 -40
rect 185 -45 189 -43
rect 145 -48 160 -45
rect 156 -49 160 -48
rect 177 -48 189 -45
rect 177 -49 181 -48
rect 371 -44 375 -43
rect 286 -46 296 -45
rect 156 -52 160 -51
rect 177 -52 181 -51
rect 156 -55 159 -52
rect 286 -49 296 -48
rect 339 -49 343 -48
rect 298 -53 299 -49
rect 303 -53 304 -49
rect 314 -53 316 -49
rect 339 -52 343 -51
rect 306 -54 316 -53
rect 327 -56 396 -52
rect 306 -57 316 -56
rect 331 -57 335 -56
rect 331 -60 335 -59
rect 347 -78 351 -77
rect 37 -84 40 -82
rect 39 -95 40 -84
rect 42 -95 43 -82
rect 53 -84 56 -82
rect 35 -98 39 -97
rect 35 -103 39 -102
rect 31 -118 32 -105
rect 34 -118 35 -105
rect 55 -95 56 -84
rect 58 -95 59 -82
rect 69 -84 72 -82
rect 51 -98 55 -97
rect 51 -103 55 -102
rect 47 -118 48 -105
rect 50 -118 51 -105
rect 71 -95 72 -84
rect 74 -95 75 -82
rect 85 -84 88 -82
rect 67 -98 71 -97
rect 67 -103 71 -102
rect 63 -118 64 -105
rect 66 -118 67 -105
rect 87 -95 88 -84
rect 90 -95 91 -82
rect 101 -84 104 -82
rect 83 -98 87 -97
rect 83 -103 87 -102
rect 79 -118 80 -105
rect 82 -118 83 -105
rect 103 -95 104 -84
rect 106 -95 107 -82
rect 340 -92 344 -80
rect 346 -87 347 -80
rect 363 -78 367 -77
rect 346 -92 350 -87
rect 340 -95 343 -92
rect 99 -98 103 -97
rect 99 -103 103 -102
rect 95 -118 96 -105
rect 98 -118 99 -105
rect 332 -97 336 -95
rect 335 -105 336 -97
rect 338 -105 343 -95
rect 356 -92 360 -80
rect 362 -87 363 -80
rect 379 -78 383 -77
rect 362 -92 366 -87
rect 356 -95 359 -92
rect 348 -97 352 -95
rect 351 -105 352 -97
rect 354 -105 359 -95
rect 372 -92 376 -80
rect 378 -87 379 -80
rect 395 -78 399 -77
rect 378 -92 382 -87
rect 372 -95 375 -92
rect 364 -97 368 -95
rect 367 -105 368 -97
rect 370 -105 375 -95
rect 335 -257 336 -247
rect 332 -259 336 -257
rect 338 -259 343 -247
rect 47 -267 48 -263
rect 41 -268 45 -267
rect 63 -267 64 -263
rect 57 -268 61 -267
rect 79 -267 80 -263
rect 73 -268 77 -267
rect 95 -267 96 -263
rect 89 -268 93 -267
rect 111 -267 112 -263
rect 340 -262 343 -259
rect 388 -92 392 -80
rect 394 -87 395 -80
rect 394 -92 398 -87
rect 388 -95 391 -92
rect 380 -97 384 -95
rect 383 -105 384 -97
rect 386 -105 391 -95
rect 351 -257 352 -247
rect 348 -259 352 -257
rect 354 -259 359 -247
rect 105 -268 109 -267
rect 41 -273 45 -270
rect 57 -273 61 -270
rect 73 -273 77 -270
rect 89 -273 93 -270
rect 105 -273 109 -270
rect 41 -276 45 -275
rect 41 -279 42 -276
rect 57 -276 61 -275
rect 57 -279 58 -276
rect 73 -276 77 -275
rect 73 -279 74 -276
rect 89 -276 93 -275
rect 89 -279 90 -276
rect 340 -274 344 -262
rect 346 -267 350 -262
rect 356 -262 359 -259
rect 367 -257 368 -247
rect 364 -259 368 -257
rect 370 -259 375 -247
rect 346 -274 347 -267
rect 105 -276 109 -275
rect 356 -274 360 -262
rect 362 -267 366 -262
rect 372 -262 375 -259
rect 383 -257 384 -247
rect 380 -259 384 -257
rect 386 -259 391 -247
rect 362 -274 363 -267
rect 372 -274 376 -262
rect 378 -267 382 -262
rect 388 -262 391 -259
rect 378 -274 379 -267
rect 388 -274 392 -262
rect 394 -267 398 -262
rect 394 -274 395 -267
rect 105 -279 106 -276
rect 347 -277 351 -276
rect 363 -277 367 -276
rect 379 -277 383 -276
rect 395 -277 399 -276
<< pdiffusion >>
rect 329 28 393 29
rect 331 23 335 24
rect 339 23 343 24
rect 347 23 351 24
rect 355 23 359 24
rect 363 23 367 24
rect 371 23 375 24
rect 379 23 383 24
rect 387 23 391 24
rect 331 20 335 21
rect 339 20 343 21
rect 347 20 351 21
rect 355 20 359 21
rect 363 20 367 21
rect 371 20 375 21
rect 379 20 383 21
rect 387 20 391 21
rect 126 8 127 12
rect 4 -64 5 0
rect 9 -6 10 -2
rect 12 -6 13 -2
rect 9 -14 10 -10
rect 12 -14 13 -10
rect 9 -22 10 -18
rect 12 -22 13 -18
rect 9 -30 10 -26
rect 12 -30 13 -26
rect 9 -38 10 -34
rect 12 -38 13 -34
rect 9 -46 10 -42
rect 12 -46 13 -42
rect 9 -54 10 -50
rect 12 -54 13 -50
rect 9 -62 10 -58
rect 12 -62 13 -58
rect 129 7 133 8
rect 129 4 133 5
rect 207 8 208 12
rect 201 7 205 8
rect 129 -1 133 0
rect 201 4 205 5
rect 254 3 259 7
rect 201 -1 205 0
rect 254 2 274 3
rect 254 -1 274 0
rect 129 -4 133 -3
rect 201 -4 205 -3
rect 126 -8 127 -4
rect 129 -9 133 -8
rect 129 -12 133 -11
rect 207 -8 208 -4
rect 224 -5 226 -1
rect 246 -5 247 -1
rect 251 -5 252 -1
rect 201 -9 205 -8
rect 224 -6 244 -5
rect 224 -9 244 -8
rect 129 -17 133 -16
rect 201 -12 205 -11
rect 224 -13 226 -9
rect 254 -13 259 -9
rect 201 -17 205 -16
rect 254 -14 274 -13
rect 254 -17 274 -16
rect 129 -20 133 -19
rect 201 -20 205 -19
rect 126 -24 127 -20
rect 129 -25 133 -24
rect 129 -28 133 -27
rect 207 -24 208 -20
rect 224 -21 226 -17
rect 246 -21 247 -17
rect 251 -21 252 -17
rect 201 -25 205 -24
rect 224 -22 244 -21
rect 224 -25 244 -24
rect 129 -33 133 -32
rect 201 -28 205 -27
rect 224 -29 226 -25
rect 254 -29 259 -25
rect 201 -33 205 -32
rect 254 -30 274 -29
rect 254 -33 274 -32
rect 129 -36 133 -35
rect 201 -36 205 -35
rect 126 -40 127 -36
rect 129 -41 133 -40
rect 129 -44 133 -43
rect 207 -40 208 -36
rect 224 -37 226 -33
rect 246 -37 247 -33
rect 251 -37 252 -33
rect 201 -41 205 -40
rect 224 -38 244 -37
rect 224 -41 244 -40
rect 129 -49 133 -48
rect 201 -44 205 -43
rect 224 -45 226 -41
rect 254 -45 259 -41
rect 201 -49 205 -48
rect 254 -46 274 -45
rect 254 -49 274 -48
rect 129 -52 133 -51
rect 126 -56 127 -52
rect 201 -52 205 -51
rect 207 -56 208 -52
rect 224 -53 226 -49
rect 246 -53 247 -49
rect 251 -53 252 -49
rect 224 -54 244 -53
rect 224 -57 244 -56
rect 224 -61 226 -57
rect 31 -148 32 -130
rect 29 -155 32 -148
rect 34 -155 35 -130
rect 35 -158 39 -157
rect 35 -163 39 -162
rect 47 -148 48 -130
rect 45 -155 48 -148
rect 50 -155 51 -130
rect 39 -189 40 -165
rect 35 -191 40 -189
rect 42 -182 43 -165
rect 42 -191 45 -182
rect 51 -158 55 -157
rect 51 -163 55 -162
rect 63 -148 64 -130
rect 61 -155 64 -148
rect 66 -155 67 -130
rect 55 -189 56 -165
rect 51 -191 56 -189
rect 58 -182 59 -165
rect 58 -191 61 -182
rect 67 -158 71 -157
rect 67 -163 71 -162
rect 79 -148 80 -130
rect 77 -155 80 -148
rect 82 -155 83 -130
rect 71 -189 72 -165
rect 67 -191 72 -189
rect 74 -182 75 -165
rect 74 -191 77 -182
rect 83 -158 87 -157
rect 83 -163 87 -162
rect 95 -148 96 -130
rect 93 -155 96 -148
rect 98 -155 99 -130
rect 87 -189 88 -165
rect 83 -191 88 -189
rect 90 -182 91 -165
rect 90 -191 93 -182
rect 99 -158 103 -157
rect 99 -163 103 -162
rect 335 -139 336 -117
rect 332 -141 336 -139
rect 338 -141 343 -117
rect 340 -144 343 -141
rect 351 -139 352 -117
rect 348 -141 352 -139
rect 354 -141 359 -117
rect 103 -189 104 -165
rect 99 -191 104 -189
rect 106 -182 107 -165
rect 106 -191 109 -182
rect 41 -206 42 -204
rect 41 -207 45 -206
rect 57 -206 58 -204
rect 57 -207 61 -206
rect 73 -206 74 -204
rect 73 -207 77 -206
rect 89 -206 90 -204
rect 89 -207 93 -206
rect 105 -206 106 -204
rect 105 -207 109 -206
rect 41 -212 45 -209
rect 57 -212 61 -209
rect 73 -212 77 -209
rect 89 -212 93 -209
rect 105 -212 109 -209
rect 340 -168 344 -144
rect 346 -149 350 -144
rect 356 -144 359 -141
rect 367 -139 368 -117
rect 364 -141 368 -139
rect 370 -141 375 -117
rect 346 -168 347 -149
rect 347 -171 351 -170
rect 340 -209 344 -185
rect 346 -209 347 -185
rect 340 -213 343 -209
rect 41 -215 45 -214
rect 47 -219 48 -215
rect 57 -215 61 -214
rect 63 -219 64 -215
rect 73 -215 77 -214
rect 79 -219 80 -215
rect 89 -215 93 -214
rect 95 -219 96 -215
rect 105 -215 109 -214
rect 111 -219 112 -215
rect 41 -238 42 -236
rect 41 -239 45 -238
rect 57 -238 58 -236
rect 57 -239 61 -238
rect 73 -238 74 -236
rect 73 -239 77 -238
rect 89 -238 90 -236
rect 89 -239 93 -238
rect 105 -238 106 -236
rect 335 -235 336 -213
rect 338 -235 343 -213
rect 105 -239 109 -238
rect 41 -244 45 -241
rect 57 -244 61 -241
rect 73 -244 77 -241
rect 89 -244 93 -241
rect 105 -244 109 -241
rect 41 -247 45 -246
rect 47 -251 48 -247
rect 57 -247 61 -246
rect 63 -251 64 -247
rect 73 -247 77 -246
rect 79 -251 80 -247
rect 89 -247 93 -246
rect 95 -251 96 -247
rect 105 -247 109 -246
rect 111 -251 112 -247
rect 356 -168 360 -144
rect 362 -149 366 -144
rect 372 -144 375 -141
rect 383 -139 384 -117
rect 380 -141 384 -139
rect 386 -141 391 -117
rect 362 -168 363 -149
rect 363 -171 367 -170
rect 356 -209 360 -185
rect 362 -209 363 -185
rect 356 -213 359 -209
rect 351 -235 352 -213
rect 354 -235 359 -213
rect 372 -168 376 -144
rect 378 -149 382 -144
rect 388 -144 391 -141
rect 378 -168 379 -149
rect 379 -171 383 -170
rect 372 -209 376 -185
rect 378 -209 379 -185
rect 372 -213 375 -209
rect 367 -235 368 -213
rect 370 -235 375 -213
rect 388 -168 392 -144
rect 394 -149 398 -144
rect 394 -168 395 -149
rect 395 -171 399 -170
rect 388 -209 392 -185
rect 394 -209 395 -185
rect 388 -213 391 -209
rect 383 -235 384 -213
rect 386 -235 391 -213
<< metal1 >>
rect 16 26 29 30
rect 113 26 303 32
rect 329 28 393 29
rect 16 24 113 26
rect 16 16 20 24
rect 126 8 127 12
rect 137 8 145 11
rect 153 8 156 12
rect 8 7 12 8
rect 30 2 37 5
rect 41 2 53 5
rect 57 2 69 5
rect 73 2 85 5
rect 89 2 101 5
rect 105 2 109 5
rect 4 -64 5 0
rect 17 -6 93 -3
rect 97 -6 109 -3
rect 113 -6 114 -2
rect 122 -4 126 8
rect 137 4 140 8
rect 133 1 136 4
rect 126 -8 127 -4
rect 137 -8 145 -5
rect 153 -8 156 4
rect 17 -14 93 -11
rect 113 -11 115 -10
rect 97 -13 115 -11
rect 97 -14 116 -13
rect 17 -22 93 -19
rect 113 -19 114 -18
rect 97 -22 114 -19
rect 122 -20 126 -8
rect 137 -12 140 -8
rect 133 -15 136 -12
rect 126 -24 127 -20
rect 137 -24 145 -21
rect 153 -24 156 -12
rect 17 -30 77 -27
rect 81 -30 109 -27
rect 113 -29 115 -26
rect 113 -30 116 -29
rect 17 -38 77 -35
rect 113 -35 114 -34
rect 81 -38 114 -35
rect 122 -36 126 -24
rect 137 -28 140 -24
rect 133 -31 136 -28
rect 126 -40 127 -36
rect 137 -40 145 -37
rect 153 -40 156 -28
rect 17 -46 77 -43
rect 113 -43 115 -42
rect 81 -45 115 -43
rect 81 -46 116 -45
rect 17 -54 45 -51
rect 49 -54 61 -51
rect 113 -51 114 -50
rect 65 -54 114 -51
rect 122 -52 126 -40
rect 137 -44 140 -40
rect 133 -47 136 -44
rect 126 -56 127 -52
rect 17 -62 45 -59
rect 113 -59 115 -58
rect 49 -61 115 -59
rect 49 -62 116 -61
rect 122 -64 126 -56
rect 1 -185 5 -64
rect 30 -69 37 -66
rect 41 -69 53 -66
rect 57 -69 69 -66
rect 73 -69 85 -66
rect 89 -69 101 -66
rect 105 -69 119 -66
rect 122 -68 131 -64
rect 8 -72 12 -71
rect 116 -76 119 -69
rect 1 -215 5 -189
rect 9 -207 12 -76
rect 35 -77 39 -76
rect 43 -77 47 -76
rect 51 -77 55 -76
rect 59 -77 63 -76
rect 67 -77 71 -76
rect 75 -77 79 -76
rect 83 -77 87 -76
rect 91 -77 95 -76
rect 99 -77 103 -76
rect 107 -77 111 -76
rect 43 -82 47 -81
rect 59 -82 63 -81
rect 35 -98 39 -97
rect 75 -82 79 -81
rect 51 -98 55 -97
rect 91 -82 95 -81
rect 67 -98 71 -97
rect 107 -82 111 -81
rect 83 -98 87 -97
rect 123 -84 131 -68
rect 153 -68 156 -44
rect 163 -76 167 26
rect 170 -4 174 -3
rect 177 -4 181 26
rect 208 15 292 19
rect 208 12 212 15
rect 189 8 195 11
rect 207 8 208 12
rect 192 4 195 8
rect 196 1 201 4
rect 208 -4 212 8
rect 252 -1 256 15
rect 299 10 303 26
rect 326 24 329 28
rect 393 24 395 28
rect 318 17 322 20
rect 398 20 402 21
rect 274 4 286 7
rect 277 -1 280 4
rect 299 6 322 10
rect 299 -1 303 6
rect 189 -8 195 -5
rect 207 -8 208 -4
rect 246 -5 247 -1
rect 251 -5 252 -1
rect 298 -5 299 -1
rect 303 -5 304 -1
rect 321 -5 322 -1
rect 170 -20 174 -19
rect 177 -20 181 -8
rect 192 -12 195 -8
rect 196 -15 201 -12
rect 208 -20 212 -8
rect 244 -13 245 -9
rect 252 -17 256 -5
rect 274 -12 286 -9
rect 277 -17 280 -12
rect 299 -17 303 -5
rect 316 -13 317 -9
rect 321 -13 322 -9
rect 189 -24 195 -21
rect 207 -24 208 -20
rect 246 -21 247 -17
rect 251 -21 252 -17
rect 298 -21 299 -17
rect 303 -21 304 -17
rect 321 -21 322 -17
rect 170 -36 174 -35
rect 177 -36 181 -24
rect 192 -28 195 -24
rect 196 -31 201 -28
rect 208 -36 212 -24
rect 244 -29 245 -25
rect 252 -33 256 -21
rect 274 -28 286 -25
rect 277 -33 280 -28
rect 299 -33 303 -21
rect 316 -29 317 -25
rect 321 -29 322 -25
rect 189 -40 195 -37
rect 207 -40 208 -36
rect 246 -37 247 -33
rect 251 -37 252 -33
rect 298 -37 299 -33
rect 303 -37 304 -33
rect 321 -37 322 -33
rect 170 -52 174 -51
rect 177 -52 181 -40
rect 192 -44 195 -40
rect 196 -47 201 -44
rect 208 -52 212 -40
rect 244 -45 245 -41
rect 252 -49 256 -37
rect 274 -44 286 -41
rect 277 -49 280 -44
rect 299 -49 303 -37
rect 316 -45 317 -41
rect 321 -45 322 -41
rect 207 -56 208 -52
rect 246 -53 247 -49
rect 251 -53 252 -49
rect 298 -53 299 -49
rect 303 -53 304 -49
rect 321 -53 322 -49
rect 123 -88 127 -84
rect 99 -98 103 -97
rect 9 -239 12 -211
rect 20 -102 35 -98
rect 39 -102 51 -98
rect 55 -102 67 -98
rect 71 -102 83 -98
rect 87 -102 99 -98
rect 103 -102 116 -98
rect 16 -263 20 -102
rect 35 -103 39 -102
rect 51 -103 55 -102
rect 67 -103 71 -102
rect 83 -103 87 -102
rect 99 -103 103 -102
rect 27 -123 30 -118
rect 27 -126 35 -123
rect 43 -123 46 -118
rect 43 -126 51 -123
rect 59 -123 62 -118
rect 59 -126 67 -123
rect 75 -123 78 -118
rect 75 -126 83 -123
rect 91 -123 94 -118
rect 91 -126 99 -123
rect 27 -130 30 -126
rect 43 -130 46 -126
rect 59 -130 62 -126
rect 75 -130 78 -126
rect 91 -130 94 -126
rect 107 -130 110 -118
rect 29 -155 35 -151
rect 39 -155 51 -151
rect 35 -158 39 -157
rect 55 -155 67 -151
rect 51 -158 55 -157
rect 71 -155 83 -151
rect 67 -158 71 -157
rect 87 -155 99 -151
rect 83 -158 87 -157
rect 123 -151 131 -88
rect 103 -155 131 -151
rect 99 -158 103 -157
rect 35 -163 39 -162
rect 29 -189 35 -185
rect 43 -163 47 -162
rect 51 -163 55 -162
rect 39 -189 51 -185
rect 59 -163 63 -162
rect 67 -163 71 -162
rect 55 -189 67 -185
rect 75 -163 79 -162
rect 83 -163 87 -162
rect 71 -189 83 -185
rect 91 -163 95 -162
rect 99 -163 103 -162
rect 87 -189 99 -185
rect 107 -163 111 -162
rect 123 -185 131 -155
rect 103 -189 127 -185
rect 33 -197 37 -196
rect 41 -197 45 -196
rect 49 -197 53 -196
rect 57 -197 61 -196
rect 65 -197 69 -196
rect 73 -197 77 -196
rect 81 -197 85 -196
rect 89 -197 93 -196
rect 97 -197 101 -196
rect 105 -197 109 -196
rect 42 -202 45 -201
rect 58 -202 61 -201
rect 74 -202 77 -201
rect 90 -202 93 -201
rect 106 -202 109 -201
rect 35 -209 39 -208
rect 51 -209 55 -208
rect 67 -209 71 -208
rect 83 -209 87 -208
rect 99 -209 103 -208
rect 29 -211 116 -209
rect 26 -212 116 -211
rect 123 -215 131 -189
rect 29 -219 32 -215
rect 36 -219 41 -215
rect 47 -219 48 -215
rect 52 -219 57 -215
rect 63 -219 64 -215
rect 68 -219 73 -215
rect 79 -219 80 -215
rect 84 -219 89 -215
rect 95 -219 96 -215
rect 100 -219 105 -215
rect 111 -219 112 -215
rect 116 -219 131 -215
rect 41 -226 42 -222
rect 57 -226 58 -222
rect 73 -226 74 -222
rect 89 -226 90 -222
rect 105 -226 106 -222
rect 38 -233 45 -230
rect 54 -233 61 -230
rect 70 -233 77 -230
rect 86 -233 93 -230
rect 102 -233 109 -230
rect 42 -234 45 -233
rect 58 -234 61 -233
rect 74 -234 77 -233
rect 90 -234 93 -233
rect 106 -234 109 -233
rect 35 -241 39 -240
rect 51 -241 55 -240
rect 67 -241 71 -240
rect 83 -241 87 -240
rect 99 -241 103 -240
rect 29 -243 116 -241
rect 26 -244 116 -243
rect 123 -247 131 -219
rect 29 -251 32 -247
rect 36 -251 41 -247
rect 47 -251 48 -247
rect 52 -251 57 -247
rect 63 -251 64 -247
rect 68 -251 73 -247
rect 79 -251 80 -247
rect 84 -251 89 -247
rect 95 -251 96 -247
rect 100 -251 105 -247
rect 111 -251 112 -247
rect 116 -251 131 -247
rect 41 -260 42 -256
rect 57 -260 58 -256
rect 73 -260 74 -256
rect 89 -260 90 -256
rect 105 -260 106 -256
rect 16 -267 32 -263
rect 36 -267 41 -263
rect 47 -267 48 -263
rect 52 -267 57 -263
rect 63 -267 64 -263
rect 68 -267 73 -263
rect 79 -267 80 -263
rect 84 -267 89 -263
rect 95 -267 96 -263
rect 100 -267 105 -263
rect 111 -267 112 -263
rect 29 -273 116 -270
rect 35 -274 39 -273
rect 51 -274 55 -273
rect 67 -274 71 -273
rect 83 -274 87 -273
rect 99 -274 103 -273
rect 42 -281 45 -280
rect 58 -281 61 -280
rect 74 -281 77 -280
rect 90 -281 93 -280
rect 106 -281 109 -280
rect 38 -284 45 -281
rect 54 -284 61 -281
rect 70 -284 77 -281
rect 86 -284 93 -281
rect 102 -284 109 -281
rect 123 -284 131 -251
rect 177 -76 181 -56
rect 135 -270 138 -80
rect 163 -98 167 -80
rect 208 -84 212 -56
rect 244 -61 245 -57
rect 252 -84 256 -53
rect 299 -64 303 -53
rect 316 -61 317 -57
rect 321 -61 322 -57
rect 331 -60 334 16
rect 339 -44 342 16
rect 347 4 350 16
rect 299 -68 307 -64
rect 331 -66 335 -64
rect 339 -64 342 -48
rect 347 -64 350 0
rect 355 -12 358 16
rect 363 -12 366 16
rect 355 -28 358 -16
rect 355 -64 358 -32
rect 363 -64 366 -16
rect 371 -44 374 16
rect 379 -12 382 16
rect 371 -64 374 -48
rect 379 -64 382 -16
rect 387 -28 390 16
rect 396 4 400 6
rect 396 -4 400 0
rect 407 -5 408 -1
rect 396 -12 400 -8
rect 407 -13 408 -9
rect 396 -20 400 -16
rect 407 -21 408 -17
rect 396 -28 400 -24
rect 407 -29 408 -25
rect 387 -64 390 -32
rect 396 -36 400 -32
rect 407 -37 408 -33
rect 396 -44 400 -40
rect 407 -45 408 -41
rect 396 -52 400 -48
rect 407 -53 408 -49
rect 396 -60 400 -56
rect 407 -61 408 -57
rect 339 -66 343 -64
rect 347 -66 351 -64
rect 355 -66 359 -64
rect 363 -66 367 -64
rect 371 -66 375 -64
rect 379 -66 383 -64
rect 387 -66 391 -64
rect 292 -90 295 -72
rect 299 -73 307 -72
rect 299 -76 331 -73
rect 303 -77 331 -76
rect 335 -77 347 -73
rect 351 -77 363 -73
rect 367 -77 379 -73
rect 383 -77 395 -73
rect 303 -80 307 -77
rect 143 -240 146 -212
rect 135 -284 138 -274
rect 143 -284 146 -244
rect 284 -281 287 -146
rect 292 -261 295 -94
rect 292 -281 295 -265
rect 299 -277 307 -80
rect 347 -78 351 -77
rect 363 -78 367 -77
rect 379 -78 383 -77
rect 395 -78 399 -77
rect 327 -94 335 -91
rect 339 -94 351 -91
rect 355 -94 367 -91
rect 371 -94 383 -91
rect 387 -94 399 -91
rect 331 -110 334 -105
rect 347 -110 350 -105
rect 363 -110 366 -105
rect 379 -110 382 -105
rect 331 -117 334 -114
rect 347 -117 350 -114
rect 363 -117 366 -114
rect 379 -117 382 -114
rect 327 -146 335 -143
rect 339 -146 351 -143
rect 355 -146 367 -143
rect 371 -146 383 -143
rect 387 -146 399 -143
rect 347 -171 351 -170
rect 363 -171 367 -170
rect 379 -171 383 -170
rect 395 -171 399 -170
rect 323 -175 331 -171
rect 335 -175 347 -171
rect 351 -175 363 -171
rect 367 -175 379 -171
rect 383 -175 395 -171
rect 323 -185 327 -175
rect 343 -182 344 -178
rect 359 -182 360 -178
rect 375 -182 376 -178
rect 391 -182 392 -178
rect 327 -189 347 -185
rect 351 -189 363 -185
rect 367 -189 379 -185
rect 383 -189 395 -185
rect 331 -240 334 -235
rect 347 -240 350 -235
rect 363 -240 366 -235
rect 379 -240 382 -235
rect 331 -247 334 -244
rect 347 -247 350 -244
rect 363 -247 366 -244
rect 379 -247 382 -244
rect 327 -264 335 -261
rect 339 -264 351 -261
rect 355 -264 367 -261
rect 371 -264 383 -261
rect 387 -264 399 -261
rect 347 -277 351 -276
rect 363 -277 367 -276
rect 379 -277 383 -276
rect 395 -277 399 -276
rect 299 -281 331 -277
rect 335 -281 347 -277
rect 351 -281 363 -277
rect 367 -281 379 -277
rect 383 -281 395 -277
<< metal2 >>
rect 113 23 280 25
rect 9 22 280 23
rect 9 20 117 22
rect 9 12 12 20
rect 9 -72 12 8
rect 16 -98 20 12
rect 26 -65 29 1
rect 34 -70 37 12
rect 42 -70 45 12
rect 50 -70 53 12
rect 58 -70 61 12
rect 66 -70 69 12
rect 74 -70 77 12
rect 82 -70 85 12
rect 90 -70 93 12
rect 98 -70 101 12
rect 106 -70 109 12
rect 277 9 280 22
rect 292 24 322 28
rect 292 19 296 24
rect 318 17 398 20
rect 314 9 317 16
rect 277 6 317 9
rect 326 6 396 10
rect 140 0 181 3
rect 196 0 215 3
rect 118 -4 132 -3
rect 118 -6 170 -4
rect 129 -7 170 -6
rect 178 -5 181 0
rect 281 -4 317 -1
rect 321 -4 408 -1
rect 178 -8 215 -5
rect 140 -16 181 -13
rect 249 -13 317 -10
rect 321 -12 408 -9
rect 196 -16 215 -13
rect 118 -20 132 -19
rect 118 -22 170 -20
rect 129 -23 170 -22
rect 178 -21 181 -16
rect 281 -20 317 -17
rect 321 -20 408 -17
rect 178 -24 215 -21
rect 140 -32 181 -29
rect 249 -29 317 -26
rect 321 -28 408 -25
rect 196 -32 215 -29
rect 118 -36 132 -35
rect 118 -38 170 -36
rect 129 -39 170 -38
rect 178 -37 181 -32
rect 281 -36 317 -33
rect 321 -36 408 -33
rect 178 -40 215 -37
rect 140 -48 181 -45
rect 249 -45 317 -42
rect 321 -44 408 -41
rect 196 -48 215 -45
rect 118 -52 132 -51
rect 118 -54 170 -52
rect 129 -55 170 -54
rect 178 -53 181 -48
rect 281 -52 317 -49
rect 321 -52 408 -49
rect 178 -56 215 -53
rect 249 -61 317 -58
rect 321 -60 408 -57
rect 34 -73 38 -70
rect 42 -73 46 -70
rect 50 -73 54 -70
rect 58 -73 62 -70
rect 66 -73 70 -70
rect 74 -73 78 -70
rect 82 -73 86 -70
rect 90 -73 94 -70
rect 98 -73 102 -70
rect 106 -73 110 -70
rect 157 -72 292 -69
rect 35 -77 38 -73
rect 43 -77 46 -73
rect 51 -77 54 -73
rect 59 -77 62 -73
rect 67 -77 70 -73
rect 75 -77 78 -73
rect 83 -77 86 -73
rect 91 -77 94 -73
rect 99 -77 102 -73
rect 107 -77 110 -73
rect 120 -80 135 -77
rect 167 -80 177 -76
rect 181 -80 299 -76
rect 35 -122 38 -81
rect 43 -158 46 -81
rect 51 -122 54 -81
rect 59 -158 62 -81
rect 67 -122 70 -81
rect 75 -158 78 -81
rect 83 -122 86 -81
rect 91 -158 94 -81
rect 99 -122 102 -81
rect 107 -158 110 -81
rect 131 -88 208 -84
rect 212 -88 252 -84
rect 296 -94 323 -91
rect 120 -102 163 -98
rect 331 -103 334 -70
rect 347 -103 350 -70
rect 363 -103 366 -70
rect 379 -103 382 -70
rect 331 -106 343 -103
rect 347 -106 359 -103
rect 363 -106 375 -103
rect 379 -106 391 -103
rect 288 -146 323 -143
rect 43 -180 46 -162
rect 59 -180 62 -162
rect 75 -180 78 -162
rect 91 -180 94 -162
rect 107 -180 110 -162
rect 34 -183 46 -180
rect 50 -183 62 -180
rect 66 -183 78 -180
rect 82 -183 94 -180
rect 98 -183 110 -180
rect 5 -189 25 -185
rect 34 -197 37 -183
rect 50 -197 53 -183
rect 66 -197 69 -183
rect 82 -197 85 -183
rect 98 -197 101 -183
rect 131 -189 323 -185
rect 41 -205 44 -201
rect 57 -205 60 -201
rect 73 -205 76 -201
rect 89 -205 92 -201
rect 105 -205 108 -201
rect 12 -211 25 -208
rect 34 -208 44 -205
rect 50 -208 60 -205
rect 66 -208 76 -205
rect 82 -208 92 -205
rect 98 -208 108 -205
rect 5 -219 25 -215
rect 34 -229 37 -208
rect 12 -243 25 -240
rect 34 -281 37 -233
rect 42 -256 45 -226
rect 50 -229 53 -208
rect 42 -284 45 -260
rect 50 -281 53 -233
rect 58 -256 61 -226
rect 66 -229 69 -208
rect 58 -284 61 -260
rect 66 -281 69 -233
rect 74 -256 77 -226
rect 82 -229 85 -208
rect 74 -284 77 -260
rect 82 -281 85 -233
rect 90 -256 93 -226
rect 98 -229 101 -208
rect 120 -212 142 -209
rect 331 -213 334 -114
rect 340 -178 343 -106
rect 347 -213 350 -114
rect 356 -178 359 -106
rect 363 -213 366 -114
rect 372 -178 375 -106
rect 379 -213 382 -114
rect 388 -178 391 -106
rect 331 -216 342 -213
rect 347 -216 358 -213
rect 363 -216 374 -213
rect 379 -216 390 -213
rect 90 -284 93 -260
rect 98 -281 101 -233
rect 106 -256 109 -226
rect 120 -244 142 -241
rect 106 -284 109 -260
rect 296 -264 323 -261
rect 120 -273 135 -270
rect 331 -281 334 -244
rect 339 -281 342 -216
rect 347 -281 350 -244
rect 355 -281 358 -216
rect 363 -281 366 -244
rect 371 -281 374 -216
rect 379 -281 382 -244
rect 387 -281 390 -216
<< ntransistor >>
rect 42 -54 44 -50
rect 42 -62 44 -58
rect 50 -62 52 -58
rect 66 -54 68 -50
rect 90 -6 92 -2
rect 145 5 149 7
rect 185 5 189 7
rect 106 -6 108 -2
rect 156 -3 160 -1
rect 286 0 296 2
rect 177 -3 181 -1
rect 90 -14 92 -10
rect 98 -14 100 -10
rect 82 -30 84 -26
rect 82 -38 84 -34
rect 82 -46 84 -42
rect 98 -22 100 -18
rect 145 -11 149 -9
rect 347 -3 351 -1
rect 306 -8 316 -6
rect 185 -11 189 -9
rect 156 -19 160 -17
rect 355 -11 359 -9
rect 363 -11 367 -9
rect 286 -16 296 -14
rect 177 -19 181 -17
rect 106 -30 108 -26
rect 145 -27 149 -25
rect 379 -19 383 -17
rect 306 -24 316 -22
rect 185 -27 189 -25
rect 156 -35 160 -33
rect 387 -27 391 -25
rect 286 -32 296 -30
rect 177 -35 181 -33
rect 145 -43 149 -41
rect 355 -35 359 -33
rect 306 -40 316 -38
rect 185 -43 189 -41
rect 156 -51 160 -49
rect 371 -43 375 -41
rect 286 -48 296 -46
rect 177 -51 181 -49
rect 339 -51 343 -49
rect 306 -56 316 -54
rect 331 -59 335 -57
rect 40 -95 42 -82
rect 32 -118 34 -105
rect 56 -95 58 -82
rect 48 -118 50 -105
rect 72 -95 74 -82
rect 64 -118 66 -105
rect 88 -95 90 -82
rect 80 -118 82 -105
rect 104 -95 106 -82
rect 344 -92 346 -80
rect 96 -118 98 -105
rect 336 -105 338 -95
rect 360 -92 362 -80
rect 352 -105 354 -95
rect 376 -92 378 -80
rect 368 -105 370 -95
rect 336 -259 338 -247
rect 392 -92 394 -80
rect 384 -105 386 -95
rect 352 -259 354 -247
rect 41 -270 45 -268
rect 57 -270 61 -268
rect 73 -270 77 -268
rect 89 -270 93 -268
rect 105 -270 109 -268
rect 41 -275 45 -273
rect 57 -275 61 -273
rect 73 -275 77 -273
rect 89 -275 93 -273
rect 105 -275 109 -273
rect 344 -274 346 -262
rect 368 -259 370 -247
rect 360 -274 362 -262
rect 384 -259 386 -247
rect 376 -274 378 -262
rect 392 -274 394 -262
<< ptransistor >>
rect 331 21 335 23
rect 339 21 343 23
rect 347 21 351 23
rect 355 21 359 23
rect 363 21 367 23
rect 371 21 375 23
rect 379 21 383 23
rect 387 21 391 23
rect 10 -6 12 -2
rect 10 -14 12 -10
rect 10 -22 12 -18
rect 10 -30 12 -26
rect 10 -38 12 -34
rect 10 -46 12 -42
rect 10 -54 12 -50
rect 10 -62 12 -58
rect 129 5 133 7
rect 201 5 205 7
rect 129 -3 133 -1
rect 254 0 274 2
rect 201 -3 205 -1
rect 129 -11 133 -9
rect 224 -8 244 -6
rect 201 -11 205 -9
rect 129 -19 133 -17
rect 254 -16 274 -14
rect 201 -19 205 -17
rect 129 -27 133 -25
rect 224 -24 244 -22
rect 201 -27 205 -25
rect 129 -35 133 -33
rect 254 -32 274 -30
rect 201 -35 205 -33
rect 129 -43 133 -41
rect 224 -40 244 -38
rect 201 -43 205 -41
rect 129 -51 133 -49
rect 254 -48 274 -46
rect 201 -51 205 -49
rect 224 -56 244 -54
rect 32 -155 34 -130
rect 48 -155 50 -130
rect 40 -191 42 -165
rect 64 -155 66 -130
rect 56 -191 58 -165
rect 80 -155 82 -130
rect 72 -191 74 -165
rect 96 -155 98 -130
rect 88 -191 90 -165
rect 336 -141 338 -117
rect 352 -141 354 -117
rect 104 -191 106 -165
rect 41 -209 45 -207
rect 57 -209 61 -207
rect 73 -209 77 -207
rect 89 -209 93 -207
rect 105 -209 109 -207
rect 41 -214 45 -212
rect 57 -214 61 -212
rect 73 -214 77 -212
rect 89 -214 93 -212
rect 105 -214 109 -212
rect 344 -168 346 -144
rect 368 -141 370 -117
rect 344 -209 346 -185
rect 41 -241 45 -239
rect 57 -241 61 -239
rect 73 -241 77 -239
rect 89 -241 93 -239
rect 336 -235 338 -213
rect 105 -241 109 -239
rect 41 -246 45 -244
rect 57 -246 61 -244
rect 73 -246 77 -244
rect 89 -246 93 -244
rect 105 -246 109 -244
rect 360 -168 362 -144
rect 384 -141 386 -117
rect 360 -209 362 -185
rect 352 -235 354 -213
rect 376 -168 378 -144
rect 376 -209 378 -185
rect 368 -235 370 -213
rect 392 -168 394 -144
rect 392 -209 394 -185
rect 384 -235 386 -213
<< polycontact >>
rect 398 21 402 25
rect 322 17 326 21
rect 34 8 38 12
rect 42 8 46 12
rect 50 8 54 12
rect 58 8 62 12
rect 66 8 70 12
rect 74 8 78 12
rect 82 8 86 12
rect 90 8 94 12
rect 98 8 102 12
rect 106 8 110 12
rect 8 3 12 7
rect 8 -71 12 -67
rect 152 4 156 8
rect 170 -3 174 1
rect 219 -1 223 3
rect 115 -13 119 -9
rect 152 -12 156 -8
rect 322 -5 326 -1
rect 219 -9 223 -5
rect 403 -5 407 -1
rect 170 -19 174 -15
rect 219 -17 223 -13
rect 322 -13 326 -9
rect 403 -13 407 -9
rect 115 -29 119 -25
rect 152 -28 156 -24
rect 322 -21 326 -17
rect 219 -25 223 -21
rect 403 -21 407 -17
rect 170 -35 174 -31
rect 219 -33 223 -29
rect 322 -29 326 -25
rect 403 -29 407 -25
rect 115 -45 119 -41
rect 152 -44 156 -40
rect 322 -37 326 -33
rect 219 -41 223 -37
rect 403 -37 407 -33
rect 170 -51 174 -47
rect 219 -49 223 -45
rect 322 -45 326 -41
rect 403 -45 407 -41
rect 115 -61 119 -57
rect 322 -53 326 -49
rect 219 -57 223 -53
rect 403 -53 407 -49
rect 322 -61 326 -57
rect 403 -61 407 -57
rect 339 -70 343 -66
rect 355 -70 359 -66
rect 371 -70 375 -66
rect 387 -70 391 -66
rect 34 -76 38 -72
rect 42 -76 46 -72
rect 50 -76 54 -72
rect 58 -76 62 -72
rect 66 -76 70 -72
rect 74 -76 78 -72
rect 82 -76 86 -72
rect 90 -76 94 -72
rect 98 -76 102 -72
rect 106 -76 110 -72
rect 335 -94 339 -90
rect 335 -146 339 -142
rect 351 -94 355 -90
rect 32 -196 36 -192
rect 40 -196 44 -192
rect 48 -196 52 -192
rect 56 -196 60 -192
rect 64 -196 68 -192
rect 72 -196 76 -192
rect 80 -196 84 -192
rect 88 -196 92 -192
rect 96 -196 100 -192
rect 104 -196 108 -192
rect 35 -208 39 -204
rect 51 -208 55 -204
rect 67 -208 71 -204
rect 83 -208 87 -204
rect 99 -208 103 -204
rect 351 -146 355 -142
rect 367 -94 371 -90
rect 344 -182 348 -178
rect 37 -226 41 -222
rect 53 -226 57 -222
rect 69 -226 73 -222
rect 85 -226 89 -222
rect 101 -226 105 -222
rect 35 -240 39 -236
rect 51 -240 55 -236
rect 67 -240 71 -236
rect 83 -240 87 -236
rect 99 -240 103 -236
rect 37 -260 41 -256
rect 53 -260 57 -256
rect 69 -260 73 -256
rect 85 -260 89 -256
rect 101 -260 105 -256
rect 335 -264 339 -260
rect 367 -146 371 -142
rect 383 -94 387 -90
rect 360 -182 364 -178
rect 35 -278 39 -274
rect 51 -278 55 -274
rect 67 -278 71 -274
rect 83 -278 87 -274
rect 99 -278 103 -274
rect 351 -264 355 -260
rect 383 -146 387 -142
rect 376 -182 380 -178
rect 367 -264 371 -260
rect 392 -182 396 -178
rect 383 -264 387 -260
<< ndcontact >>
rect 37 1 41 5
rect 45 -54 49 -50
rect 53 1 57 5
rect 45 -62 49 -58
rect 37 -69 41 -65
rect 53 -69 57 -65
rect 69 1 73 5
rect 61 -54 65 -50
rect 69 -69 73 -65
rect 85 1 89 5
rect 93 -6 97 -2
rect 101 1 105 5
rect 145 8 149 12
rect 185 8 189 12
rect 109 -6 113 -2
rect 286 3 296 7
rect 347 0 351 4
rect 93 -14 97 -10
rect 77 -30 81 -26
rect 77 -38 81 -34
rect 77 -46 81 -42
rect 85 -69 89 -65
rect 93 -22 97 -18
rect 145 -8 149 -4
rect 159 -8 163 -4
rect 177 -8 181 -4
rect 185 -8 189 -4
rect 286 -5 298 -1
rect 304 -5 314 -1
rect 396 -8 400 -4
rect 286 -13 296 -9
rect 306 -13 316 -9
rect 355 -16 359 -12
rect 363 -16 367 -12
rect 379 -16 383 -12
rect 109 -30 113 -26
rect 145 -24 149 -20
rect 159 -24 163 -20
rect 177 -24 181 -20
rect 185 -24 189 -20
rect 101 -69 105 -65
rect 286 -21 298 -17
rect 304 -21 314 -17
rect 396 -24 400 -20
rect 286 -29 296 -25
rect 306 -29 316 -25
rect 355 -32 359 -28
rect 387 -32 391 -28
rect 145 -40 149 -36
rect 159 -40 163 -36
rect 177 -40 181 -36
rect 185 -40 189 -36
rect 286 -37 298 -33
rect 304 -37 314 -33
rect 396 -40 400 -36
rect 286 -45 296 -41
rect 306 -45 316 -41
rect 339 -48 343 -44
rect 371 -48 375 -44
rect 159 -56 163 -52
rect 177 -56 181 -52
rect 286 -53 298 -49
rect 304 -53 314 -49
rect 396 -56 400 -52
rect 306 -61 316 -57
rect 331 -64 335 -60
rect 35 -97 39 -84
rect 43 -95 47 -82
rect 27 -118 31 -105
rect 35 -118 39 -103
rect 51 -97 55 -84
rect 59 -95 63 -82
rect 43 -118 47 -105
rect 51 -118 55 -103
rect 67 -97 71 -84
rect 75 -95 79 -82
rect 59 -118 63 -105
rect 67 -118 71 -103
rect 83 -97 87 -84
rect 91 -95 95 -82
rect 75 -118 79 -105
rect 83 -118 87 -103
rect 99 -97 103 -84
rect 107 -95 111 -82
rect 347 -87 351 -78
rect 91 -118 95 -105
rect 99 -118 103 -103
rect 331 -105 335 -97
rect 107 -118 111 -105
rect 363 -87 367 -78
rect 347 -105 351 -97
rect 379 -87 383 -78
rect 363 -105 367 -97
rect 331 -257 335 -247
rect 41 -267 47 -263
rect 57 -267 63 -263
rect 73 -267 79 -263
rect 89 -267 95 -263
rect 105 -267 111 -263
rect 395 -87 399 -78
rect 379 -105 383 -97
rect 347 -257 351 -247
rect 42 -280 46 -276
rect 58 -280 62 -276
rect 74 -280 78 -276
rect 90 -280 94 -276
rect 363 -257 367 -247
rect 347 -276 351 -267
rect 379 -257 383 -247
rect 363 -276 367 -267
rect 379 -276 383 -267
rect 395 -276 399 -267
rect 106 -280 110 -276
<< pdcontact >>
rect 329 24 393 28
rect 331 16 335 20
rect 339 16 343 20
rect 347 16 351 20
rect 355 16 359 20
rect 363 16 367 20
rect 371 16 375 20
rect 379 16 383 20
rect 387 16 391 20
rect 127 8 133 12
rect 5 -64 9 0
rect 13 -6 17 -2
rect 13 -14 17 -10
rect 13 -22 17 -18
rect 13 -30 17 -26
rect 13 -38 17 -34
rect 13 -46 17 -42
rect 13 -54 17 -50
rect 13 -62 17 -58
rect 129 0 133 4
rect 201 8 207 12
rect 201 0 205 4
rect 259 3 274 7
rect 127 -8 133 -4
rect 129 -16 133 -12
rect 201 -8 207 -4
rect 226 -5 246 -1
rect 252 -5 274 -1
rect 201 -16 205 -12
rect 226 -13 244 -9
rect 259 -13 274 -9
rect 127 -24 133 -20
rect 129 -32 133 -28
rect 201 -24 207 -20
rect 226 -21 246 -17
rect 252 -21 274 -17
rect 201 -32 205 -28
rect 226 -29 244 -25
rect 259 -29 274 -25
rect 127 -40 133 -36
rect 129 -48 133 -44
rect 201 -40 207 -36
rect 226 -37 246 -33
rect 252 -37 274 -33
rect 201 -48 205 -44
rect 226 -45 244 -41
rect 259 -45 274 -41
rect 127 -56 133 -52
rect 201 -56 207 -52
rect 226 -53 246 -49
rect 252 -53 274 -49
rect 226 -61 244 -57
rect 27 -148 31 -130
rect 35 -157 39 -130
rect 35 -189 39 -163
rect 43 -148 47 -130
rect 43 -182 47 -163
rect 51 -157 55 -130
rect 51 -189 55 -163
rect 59 -148 63 -130
rect 59 -182 63 -163
rect 67 -157 71 -130
rect 67 -189 71 -163
rect 75 -148 79 -130
rect 75 -182 79 -163
rect 83 -157 87 -130
rect 83 -189 87 -163
rect 91 -148 95 -130
rect 91 -182 95 -163
rect 99 -157 103 -130
rect 99 -189 103 -163
rect 107 -148 111 -130
rect 331 -139 335 -117
rect 347 -139 351 -117
rect 107 -182 111 -163
rect 42 -206 46 -202
rect 58 -206 62 -202
rect 74 -206 78 -202
rect 90 -206 94 -202
rect 106 -206 110 -202
rect 363 -139 367 -117
rect 347 -170 351 -149
rect 347 -209 351 -185
rect 41 -219 47 -215
rect 57 -219 63 -215
rect 73 -219 79 -215
rect 89 -219 95 -215
rect 105 -219 111 -215
rect 42 -238 46 -234
rect 58 -238 62 -234
rect 74 -238 78 -234
rect 90 -238 94 -234
rect 106 -238 110 -234
rect 331 -235 335 -213
rect 41 -251 47 -247
rect 57 -251 63 -247
rect 73 -251 79 -247
rect 89 -251 95 -247
rect 105 -251 111 -247
rect 379 -139 383 -117
rect 363 -170 367 -149
rect 363 -209 367 -185
rect 347 -235 351 -213
rect 379 -170 383 -149
rect 379 -209 383 -185
rect 363 -235 367 -213
rect 395 -170 399 -149
rect 395 -209 399 -185
rect 379 -235 383 -213
<< m2contact >>
rect 16 12 20 16
rect 34 12 38 16
rect 8 8 12 12
rect 42 12 46 16
rect 50 12 54 16
rect 58 12 62 16
rect 66 12 70 16
rect 74 12 78 16
rect 82 12 86 16
rect 90 12 94 16
rect 98 12 102 16
rect 106 12 110 16
rect 26 1 30 5
rect 114 -6 118 -2
rect 136 0 140 4
rect 114 -22 118 -18
rect 136 -16 140 -12
rect 114 -38 118 -34
rect 136 -32 140 -28
rect 114 -54 118 -50
rect 136 -48 140 -44
rect 26 -69 30 -65
rect 8 -76 12 -72
rect 1 -189 5 -185
rect 35 -81 39 -77
rect 43 -81 47 -77
rect 51 -81 55 -77
rect 59 -81 63 -77
rect 67 -81 71 -77
rect 75 -81 79 -77
rect 83 -81 87 -77
rect 91 -81 95 -77
rect 99 -81 103 -77
rect 107 -81 111 -77
rect 116 -80 120 -76
rect 153 -72 157 -68
rect 170 -8 174 -4
rect 292 15 296 19
rect 192 0 196 4
rect 215 -1 219 3
rect 322 24 326 28
rect 314 16 318 20
rect 398 16 402 20
rect 322 6 326 10
rect 277 -5 281 -1
rect 317 -5 321 -1
rect 170 -24 174 -20
rect 192 -16 196 -12
rect 215 -9 219 -5
rect 245 -13 249 -9
rect 215 -17 219 -13
rect 317 -13 321 -9
rect 277 -21 281 -17
rect 317 -21 321 -17
rect 170 -40 174 -36
rect 192 -32 196 -28
rect 215 -25 219 -21
rect 245 -29 249 -25
rect 215 -33 219 -29
rect 317 -29 321 -25
rect 277 -37 281 -33
rect 317 -37 321 -33
rect 170 -56 174 -52
rect 192 -48 196 -44
rect 215 -41 219 -37
rect 245 -45 249 -41
rect 215 -49 219 -45
rect 317 -45 321 -41
rect 277 -53 281 -49
rect 317 -53 321 -49
rect 127 -88 131 -84
rect 8 -211 12 -207
rect 1 -219 5 -215
rect 8 -243 12 -239
rect 16 -102 20 -98
rect 116 -102 120 -98
rect 35 -126 39 -122
rect 51 -126 55 -122
rect 67 -126 71 -122
rect 83 -126 87 -122
rect 99 -126 103 -122
rect 25 -189 29 -185
rect 43 -162 47 -158
rect 59 -162 63 -158
rect 75 -162 79 -158
rect 91 -162 95 -158
rect 107 -162 111 -158
rect 127 -189 131 -185
rect 33 -201 37 -197
rect 41 -201 45 -197
rect 49 -201 53 -197
rect 57 -201 61 -197
rect 65 -201 69 -197
rect 73 -201 77 -197
rect 81 -201 85 -197
rect 89 -201 93 -197
rect 97 -201 101 -197
rect 105 -201 109 -197
rect 25 -211 29 -207
rect 116 -212 120 -208
rect 25 -219 29 -215
rect 42 -226 46 -222
rect 58 -226 62 -222
rect 74 -226 78 -222
rect 90 -226 94 -222
rect 106 -226 110 -222
rect 34 -233 38 -229
rect 50 -233 54 -229
rect 66 -233 70 -229
rect 82 -233 86 -229
rect 98 -233 102 -229
rect 25 -243 29 -239
rect 116 -244 120 -240
rect 42 -260 46 -256
rect 58 -260 62 -256
rect 74 -260 78 -256
rect 90 -260 94 -256
rect 106 -260 110 -256
rect 116 -274 120 -270
rect 34 -285 38 -281
rect 50 -285 54 -281
rect 66 -285 70 -281
rect 82 -285 86 -281
rect 98 -285 102 -281
rect 135 -80 139 -76
rect 163 -80 167 -76
rect 177 -80 181 -76
rect 215 -57 219 -53
rect 245 -61 249 -57
rect 208 -88 212 -84
rect 317 -61 321 -57
rect 252 -88 256 -84
rect 292 -72 296 -68
rect 331 -70 335 -66
rect 396 6 400 10
rect 408 -5 412 -1
rect 408 -13 412 -9
rect 408 -21 412 -17
rect 408 -29 412 -25
rect 408 -37 412 -33
rect 408 -45 412 -41
rect 408 -53 412 -49
rect 408 -61 412 -57
rect 347 -70 351 -66
rect 363 -70 367 -66
rect 379 -70 383 -66
rect 163 -102 167 -98
rect 299 -80 303 -76
rect 292 -94 296 -90
rect 284 -146 288 -142
rect 142 -212 146 -208
rect 142 -244 146 -240
rect 135 -274 139 -270
rect 292 -265 296 -261
rect 323 -94 327 -90
rect 331 -114 335 -110
rect 347 -114 351 -110
rect 363 -114 367 -110
rect 379 -114 383 -110
rect 323 -146 327 -142
rect 339 -182 343 -178
rect 355 -182 359 -178
rect 371 -182 375 -178
rect 387 -182 391 -178
rect 323 -189 327 -185
rect 331 -244 335 -240
rect 347 -244 351 -240
rect 363 -244 367 -240
rect 379 -244 383 -240
rect 323 -265 327 -261
<< psubstratepcontact >>
rect 29 26 113 30
rect 396 0 400 4
rect 299 -5 303 -1
rect 396 -16 400 -12
rect 299 -21 303 -17
rect 396 -32 400 -28
rect 299 -37 303 -33
rect 396 -48 400 -44
rect 299 -53 303 -49
rect 396 -64 400 -60
rect 299 -72 307 -68
rect 331 -77 335 -73
rect 347 -77 351 -73
rect 35 -102 39 -98
rect 51 -102 55 -98
rect 67 -102 71 -98
rect 83 -102 87 -98
rect 363 -77 367 -73
rect 99 -102 103 -98
rect 379 -77 383 -73
rect 395 -77 399 -73
rect 32 -267 36 -263
rect 48 -267 52 -263
rect 64 -267 68 -263
rect 80 -267 84 -263
rect 96 -267 100 -263
rect 112 -267 116 -263
rect 331 -281 335 -277
rect 347 -281 351 -277
rect 363 -281 367 -277
rect 379 -281 383 -277
rect 395 -281 399 -277
<< nsubstratencontact >>
rect 329 29 393 33
rect 122 8 126 12
rect 0 -64 4 0
rect 208 8 212 12
rect 122 -8 126 -4
rect 208 -8 212 -4
rect 247 -5 251 -1
rect 122 -24 126 -20
rect 208 -24 212 -20
rect 247 -21 251 -17
rect 122 -40 126 -36
rect 208 -40 212 -36
rect 247 -37 251 -33
rect 122 -56 126 -52
rect 208 -56 212 -52
rect 247 -53 251 -49
rect 35 -162 39 -158
rect 51 -162 55 -158
rect 67 -162 71 -158
rect 83 -162 87 -158
rect 99 -162 103 -158
rect 331 -175 335 -171
rect 347 -175 351 -171
rect 32 -219 36 -215
rect 48 -219 52 -215
rect 64 -219 68 -215
rect 80 -219 84 -215
rect 96 -219 100 -215
rect 112 -219 116 -215
rect 32 -251 36 -247
rect 48 -251 52 -247
rect 64 -251 68 -247
rect 80 -251 84 -247
rect 96 -251 100 -247
rect 112 -251 116 -247
rect 363 -175 367 -171
rect 379 -175 383 -171
rect 395 -175 399 -171
<< labels >>
rlabel metal2 42 -262 45 -262 1 RESET
rlabel metal2 58 -262 61 -262 1 load
rlabel metal2 74 -262 77 -262 1 iter
rlabel metal2 90 -262 93 -262 1 InSt0*
rlabel metal2 106 -262 109 -262 1 InSt1*
rlabel metal1 284 -280 287 -280 1 p1-
rlabel metal1 292 -280 295 -280 1 p1
rlabel metal1 143 -283 146 -283 1 p2-
rlabel metal1 135 -283 138 -283 1 p2
rlabel metal1 123 -283 131 -283 1 Vdd!
rlabel metal1 299 -280 307 -280 1 GND!
rlabel metal1 331 -238 334 -238 1 OutSt1*
rlabel metal2 339 -238 342 -238 1 OutSt0*
rlabel metal1 347 -238 350 -238 1 ready
rlabel metal2 355 -238 358 -238 1 sreg_en
rlabel metal1 363 -238 366 -238 1 sreg_latch
rlabel metal2 371 -238 374 -238 1 add_latch
rlabel metal1 379 -238 382 -238 1 in_latch
rlabel metal2 387 -238 390 -238 1 loop_latch
<< end >>
