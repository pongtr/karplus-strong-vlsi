magic
tech scmos
timestamp 1512538665
<< polysilicon >>
rect -66 1238 -64 1240
rect -58 1238 -56 1240
rect -58 1170 -56 1172
<< metal1 >>
rect -75 1240 -71 1244
rect -95 1233 -93 1236
<< metal2 >>
rect -95 1222 -93 1226
rect -95 1127 -91 1131
rect 1799 1127 1801 1131
use sreg_left_control  sreg_left_control_0
timestamp 1512534937
transform 1 0 -99 0 1 1181
box 4 -1178 99 65
use sreg_10b  sreg_10b_0
array 0 31 56 0 0 1248
timestamp 1512379799
transform 1 0 0 0 1 3
box 0 -3 56 1245
use sreg_right  sreg_right_0
timestamp 1512379879
transform 1 0 1803 0 1 2
box -11 2 -2 1155
<< labels >>
rlabel metal2 -95 1222 -95 1226 3 GND!
rlabel metal1 -95 1233 -95 1236 3 Vdd!
rlabel metal1 -73 1242 -73 1242 1 en
rlabel polysilicon -66 1239 -64 1239 1 bp
rlabel polysilicon -58 1239 -56 1239 1 phi0
rlabel polysilicon -58 1171 -56 1171 1 phi1
rlabel metal2 -93 1127 -93 1131 3 in9
rlabel metal2 1800 1127 1800 1131 7 out9
<< end >>
