magic
tech scmos
timestamp 1512379736
use addsub_one  addsub_one_0
array 0 0 196 0 9 124
timestamp 1512379586
transform 1 0 31 0 1 38
box -27 -39 169 85
<< end >>
