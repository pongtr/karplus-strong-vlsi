magic
tech scmos
timestamp 1037203492
<< pdiffusion >>
rect 32 102 38 106
rect 42 102 48 106
rect 52 102 58 106
rect 62 102 68 106
rect 72 102 77 106
rect 32 101 77 102
rect 32 97 33 101
rect 37 97 43 101
rect 47 97 53 101
rect 57 97 63 101
rect 67 97 73 101
rect 32 96 77 97
rect 32 92 38 96
rect 42 92 48 96
rect 52 92 58 96
rect 62 92 68 96
rect 72 92 77 96
rect 32 91 77 92
rect 32 87 33 91
rect 37 87 43 91
rect 47 87 53 91
rect 57 87 63 91
rect 67 87 73 91
rect 32 86 77 87
rect 32 82 38 86
rect 42 82 48 86
rect 52 82 58 86
rect 62 82 68 86
rect 72 82 77 86
rect 32 81 77 82
rect 32 77 33 81
rect 37 77 43 81
rect 47 77 53 81
rect 57 77 63 81
rect 67 77 73 81
rect 32 76 77 77
rect 32 72 38 76
rect 42 72 48 76
rect 52 72 58 76
rect 62 72 68 76
rect 72 72 77 76
rect 32 71 77 72
rect 32 67 33 71
rect 37 67 43 71
rect 47 67 53 71
rect 57 67 63 71
rect 67 67 73 71
rect 32 66 77 67
rect 32 62 38 66
rect 42 62 48 66
rect 52 62 58 66
rect 62 62 68 66
rect 72 62 77 66
rect 32 61 77 62
rect 32 57 33 61
rect 37 57 43 61
rect 47 57 53 61
rect 57 57 63 61
rect 67 57 73 61
rect 32 56 77 57
rect 32 52 38 56
rect 42 52 48 56
rect 52 52 58 56
rect 62 52 68 56
rect 72 52 77 56
rect 32 51 77 52
rect 32 47 33 51
rect 37 47 43 51
rect 47 47 53 51
rect 57 47 63 51
rect 67 47 73 51
rect 32 46 77 47
rect 32 42 38 46
rect 42 42 48 46
rect 52 42 58 46
rect 62 42 68 46
rect 72 42 77 46
rect 32 41 77 42
rect 32 37 33 41
rect 37 37 43 41
rect 47 37 53 41
rect 57 37 63 41
rect 67 37 73 41
rect 32 36 77 37
rect 32 32 38 36
rect 42 32 48 36
rect 52 32 58 36
rect 62 32 68 36
rect 72 32 77 36
rect 32 31 77 32
rect 32 27 33 31
rect 37 27 43 31
rect 47 27 53 31
rect 57 27 63 31
rect 67 27 73 31
rect 32 26 77 27
rect 32 22 38 26
rect 42 22 48 26
rect 52 22 58 26
rect 62 22 68 26
rect 72 22 77 26
rect 32 21 77 22
rect 32 17 33 21
rect 37 17 43 21
rect 47 17 53 21
rect 57 17 63 21
rect 67 17 73 21
<< pdcontact >>
rect 38 102 42 106
rect 48 102 52 106
rect 58 102 62 106
rect 68 102 72 106
rect 33 97 37 101
rect 43 97 47 101
rect 53 97 57 101
rect 63 97 67 101
rect 73 97 77 101
rect 38 92 42 96
rect 48 92 52 96
rect 58 92 62 96
rect 68 92 72 96
rect 33 87 37 91
rect 43 87 47 91
rect 53 87 57 91
rect 63 87 67 91
rect 73 87 77 91
rect 38 82 42 86
rect 48 82 52 86
rect 58 82 62 86
rect 68 82 72 86
rect 33 77 37 81
rect 43 77 47 81
rect 53 77 57 81
rect 63 77 67 81
rect 73 77 77 81
rect 38 72 42 76
rect 48 72 52 76
rect 58 72 62 76
rect 68 72 72 76
rect 33 67 37 71
rect 43 67 47 71
rect 53 67 57 71
rect 63 67 67 71
rect 73 67 77 71
rect 38 62 42 66
rect 48 62 52 66
rect 58 62 62 66
rect 68 62 72 66
rect 33 57 37 61
rect 43 57 47 61
rect 53 57 57 61
rect 63 57 67 61
rect 73 57 77 61
rect 38 52 42 56
rect 48 52 52 56
rect 58 52 62 56
rect 68 52 72 56
rect 33 47 37 51
rect 43 47 47 51
rect 53 47 57 51
rect 63 47 67 51
rect 73 47 77 51
rect 38 42 42 46
rect 48 42 52 46
rect 58 42 62 46
rect 68 42 72 46
rect 33 37 37 41
rect 43 37 47 41
rect 53 37 57 41
rect 63 37 67 41
rect 73 37 77 41
rect 38 32 42 36
rect 48 32 52 36
rect 58 32 62 36
rect 68 32 72 36
rect 33 27 37 31
rect 43 27 47 31
rect 53 27 57 31
rect 63 27 67 31
rect 73 27 77 31
rect 38 22 42 26
rect 48 22 52 26
rect 58 22 62 26
rect 68 22 72 26
rect 33 17 37 21
rect 43 17 47 21
rect 53 17 57 21
rect 63 17 67 21
rect 73 17 77 21
<< psubstratepdiff >>
rect 7 131 103 132
rect 7 127 8 131
rect 12 127 13 131
rect 17 127 18 131
rect 22 127 23 131
rect 27 127 28 131
rect 32 127 33 131
rect 37 127 38 131
rect 42 127 43 131
rect 47 127 48 131
rect 52 127 53 131
rect 57 127 58 131
rect 62 127 63 131
rect 67 127 68 131
rect 72 127 73 131
rect 77 127 78 131
rect 82 127 83 131
rect 87 127 88 131
rect 92 127 93 131
rect 97 127 98 131
rect 102 127 103 131
rect 7 126 103 127
rect 7 122 8 126
rect 12 122 13 126
rect 7 121 13 122
rect 7 117 8 121
rect 12 117 13 121
rect 97 122 98 126
rect 102 122 103 126
rect 97 121 103 122
rect 7 116 13 117
rect 7 112 8 116
rect 12 112 13 116
rect 7 111 13 112
rect 7 107 8 111
rect 12 107 13 111
rect 7 106 13 107
rect 7 102 8 106
rect 12 102 13 106
rect 7 101 13 102
rect 7 97 8 101
rect 12 97 13 101
rect 7 96 13 97
rect 7 92 8 96
rect 12 92 13 96
rect 7 91 13 92
rect 7 87 8 91
rect 12 87 13 91
rect 7 86 13 87
rect 7 82 8 86
rect 12 82 13 86
rect 7 81 13 82
rect 7 77 8 81
rect 12 77 13 81
rect 7 76 13 77
rect 7 72 8 76
rect 12 72 13 76
rect 7 71 13 72
rect 7 67 8 71
rect 12 67 13 71
rect 7 66 13 67
rect 7 62 8 66
rect 12 62 13 66
rect 7 61 13 62
rect 7 57 8 61
rect 12 57 13 61
rect 7 56 13 57
rect 7 52 8 56
rect 12 52 13 56
rect 7 51 13 52
rect 7 47 8 51
rect 12 47 13 51
rect 7 46 13 47
rect 7 42 8 46
rect 12 42 13 46
rect 7 41 13 42
rect 7 37 8 41
rect 12 37 13 41
rect 7 36 13 37
rect 7 32 8 36
rect 12 32 13 36
rect 7 31 13 32
rect 7 27 8 31
rect 12 27 13 31
rect 7 26 13 27
rect 7 22 8 26
rect 12 22 13 26
rect 7 21 13 22
rect 7 17 8 21
rect 12 17 13 21
rect 7 16 13 17
rect 7 12 8 16
rect 12 12 13 16
rect 7 11 13 12
rect 7 7 8 11
rect 12 7 13 11
rect 7 6 13 7
rect 7 2 8 6
rect 12 2 13 6
rect 97 117 98 121
rect 102 117 103 121
rect 97 116 103 117
rect 97 112 98 116
rect 102 112 103 116
rect 97 111 103 112
rect 97 107 98 111
rect 102 107 103 111
rect 97 106 103 107
rect 97 102 98 106
rect 102 102 103 106
rect 97 101 103 102
rect 97 97 98 101
rect 102 97 103 101
rect 97 96 103 97
rect 97 92 98 96
rect 102 92 103 96
rect 97 91 103 92
rect 97 87 98 91
rect 102 87 103 91
rect 97 86 103 87
rect 97 82 98 86
rect 102 82 103 86
rect 97 81 103 82
rect 97 77 98 81
rect 102 77 103 81
rect 97 76 103 77
rect 97 72 98 76
rect 102 72 103 76
rect 97 71 103 72
rect 97 67 98 71
rect 102 67 103 71
rect 97 66 103 67
rect 97 62 98 66
rect 102 62 103 66
rect 97 61 103 62
rect 97 57 98 61
rect 102 57 103 61
rect 97 56 103 57
rect 97 52 98 56
rect 102 52 103 56
rect 97 51 103 52
rect 97 47 98 51
rect 102 47 103 51
rect 97 46 103 47
rect 97 42 98 46
rect 102 42 103 46
rect 97 41 103 42
rect 97 37 98 41
rect 102 37 103 41
rect 97 36 103 37
rect 97 32 98 36
rect 102 32 103 36
rect 97 31 103 32
rect 97 27 98 31
rect 102 27 103 31
rect 97 26 103 27
rect 97 22 98 26
rect 102 22 103 26
rect 97 21 103 22
rect 97 17 98 21
rect 102 17 103 21
rect 97 16 103 17
rect 97 12 98 16
rect 102 12 103 16
rect 97 11 103 12
rect 97 7 98 11
rect 102 7 103 11
rect 97 6 103 7
rect 7 1 13 2
rect 7 -3 8 1
rect 12 -3 13 1
rect 97 2 98 6
rect 102 2 103 6
rect 97 1 103 2
rect 97 -3 98 1
rect 102 -3 103 1
rect 7 -4 103 -3
rect 7 -8 8 -4
rect 12 -8 13 -4
rect 17 -8 18 -4
rect 22 -8 23 -4
rect 27 -8 28 -4
rect 32 -8 33 -4
rect 37 -8 38 -4
rect 42 -8 43 -4
rect 47 -8 48 -4
rect 52 -8 53 -4
rect 57 -8 58 -4
rect 62 -8 63 -4
rect 67 -8 68 -4
rect 72 -8 73 -4
rect 77 -8 78 -4
rect 82 -8 83 -4
rect 87 -8 88 -4
rect 92 -8 93 -4
rect 97 -8 98 -4
rect 102 -8 103 -4
rect 7 -9 103 -8
<< nsubstratendiff >>
rect 19 118 91 120
rect 19 114 21 118
rect 25 114 28 118
rect 32 114 33 118
rect 37 114 38 118
rect 42 114 43 118
rect 47 114 48 118
rect 52 114 53 118
rect 57 114 58 118
rect 62 114 63 118
rect 67 114 68 118
rect 72 114 73 118
rect 77 114 78 118
rect 82 114 85 118
rect 89 114 91 118
rect 19 112 91 114
rect 19 111 27 112
rect 19 107 21 111
rect 25 107 27 111
rect 19 106 27 107
rect 83 111 91 112
rect 83 107 85 111
rect 89 107 91 111
rect 83 106 91 107
rect 19 102 21 106
rect 25 102 27 106
rect 19 101 27 102
rect 19 97 21 101
rect 25 97 27 101
rect 19 96 27 97
rect 19 92 21 96
rect 25 92 27 96
rect 19 91 27 92
rect 19 87 21 91
rect 25 87 27 91
rect 19 86 27 87
rect 19 82 21 86
rect 25 82 27 86
rect 19 81 27 82
rect 19 77 21 81
rect 25 77 27 81
rect 19 76 27 77
rect 19 72 21 76
rect 25 72 27 76
rect 19 71 27 72
rect 19 67 21 71
rect 25 67 27 71
rect 19 66 27 67
rect 19 62 21 66
rect 25 62 27 66
rect 19 61 27 62
rect 19 57 21 61
rect 25 57 27 61
rect 19 56 27 57
rect 19 52 21 56
rect 25 52 27 56
rect 19 51 27 52
rect 19 47 21 51
rect 25 47 27 51
rect 19 46 27 47
rect 19 42 21 46
rect 25 42 27 46
rect 19 41 27 42
rect 19 37 21 41
rect 25 37 27 41
rect 19 36 27 37
rect 19 32 21 36
rect 25 32 27 36
rect 19 31 27 32
rect 19 27 21 31
rect 25 27 27 31
rect 19 26 27 27
rect 19 22 21 26
rect 25 22 27 26
rect 19 21 27 22
rect 19 17 21 21
rect 25 17 27 21
rect 83 102 85 106
rect 89 102 91 106
rect 83 101 91 102
rect 83 97 85 101
rect 89 97 91 101
rect 83 96 91 97
rect 83 92 85 96
rect 89 92 91 96
rect 83 91 91 92
rect 83 87 85 91
rect 89 87 91 91
rect 83 86 91 87
rect 83 82 85 86
rect 89 82 91 86
rect 83 81 91 82
rect 83 77 85 81
rect 89 77 91 81
rect 83 76 91 77
rect 83 72 85 76
rect 89 72 91 76
rect 83 71 91 72
rect 83 67 85 71
rect 89 67 91 71
rect 83 66 91 67
rect 83 62 85 66
rect 89 62 91 66
rect 83 61 91 62
rect 83 57 85 61
rect 89 57 91 61
rect 83 56 91 57
rect 83 52 85 56
rect 89 52 91 56
rect 83 51 91 52
rect 83 47 85 51
rect 89 47 91 51
rect 83 46 91 47
rect 83 42 85 46
rect 89 42 91 46
rect 83 41 91 42
rect 83 37 85 41
rect 89 37 91 41
rect 83 36 91 37
rect 83 32 85 36
rect 89 32 91 36
rect 83 31 91 32
rect 83 27 85 31
rect 89 27 91 31
rect 83 26 91 27
rect 83 22 85 26
rect 89 22 91 26
rect 83 21 91 22
rect 83 17 85 21
rect 89 17 91 21
rect 19 16 27 17
rect 19 12 21 16
rect 25 12 27 16
rect 19 11 27 12
rect 83 16 91 17
rect 83 12 85 16
rect 89 12 91 16
rect 83 11 91 12
rect 19 9 91 11
rect 19 5 21 9
rect 25 5 28 9
rect 32 5 33 9
rect 37 5 38 9
rect 42 5 43 9
rect 47 5 48 9
rect 52 5 53 9
rect 57 5 58 9
rect 62 5 63 9
rect 67 5 68 9
rect 72 5 73 9
rect 77 5 78 9
rect 82 5 85 9
rect 89 5 91 9
rect 19 3 91 5
<< psubstratepcontact >>
rect 8 127 12 131
rect 13 127 17 131
rect 18 127 22 131
rect 23 127 27 131
rect 28 127 32 131
rect 33 127 37 131
rect 38 127 42 131
rect 43 127 47 131
rect 48 127 52 131
rect 53 127 57 131
rect 58 127 62 131
rect 63 127 67 131
rect 68 127 72 131
rect 73 127 77 131
rect 78 127 82 131
rect 83 127 87 131
rect 88 127 92 131
rect 93 127 97 131
rect 98 127 102 131
rect 8 122 12 126
rect 8 117 12 121
rect 98 122 102 126
rect 8 112 12 116
rect 8 107 12 111
rect 8 102 12 106
rect 8 97 12 101
rect 8 92 12 96
rect 8 87 12 91
rect 8 82 12 86
rect 8 77 12 81
rect 8 72 12 76
rect 8 67 12 71
rect 8 62 12 66
rect 8 57 12 61
rect 8 52 12 56
rect 8 47 12 51
rect 8 42 12 46
rect 8 37 12 41
rect 8 32 12 36
rect 8 27 12 31
rect 8 22 12 26
rect 8 17 12 21
rect 8 12 12 16
rect 8 7 12 11
rect 8 2 12 6
rect 98 117 102 121
rect 98 112 102 116
rect 98 107 102 111
rect 98 102 102 106
rect 98 97 102 101
rect 98 92 102 96
rect 98 87 102 91
rect 98 82 102 86
rect 98 77 102 81
rect 98 72 102 76
rect 98 67 102 71
rect 98 62 102 66
rect 98 57 102 61
rect 98 52 102 56
rect 98 47 102 51
rect 98 42 102 46
rect 98 37 102 41
rect 98 32 102 36
rect 98 27 102 31
rect 98 22 102 26
rect 98 17 102 21
rect 98 12 102 16
rect 98 7 102 11
rect 8 -3 12 1
rect 98 2 102 6
rect 98 -3 102 1
rect 8 -8 12 -4
rect 13 -8 17 -4
rect 18 -8 22 -4
rect 23 -8 27 -4
rect 28 -8 32 -4
rect 33 -8 37 -4
rect 38 -8 42 -4
rect 43 -8 47 -4
rect 48 -8 52 -4
rect 53 -8 57 -4
rect 58 -8 62 -4
rect 63 -8 67 -4
rect 68 -8 72 -4
rect 73 -8 77 -4
rect 78 -8 82 -4
rect 83 -8 87 -4
rect 88 -8 92 -4
rect 93 -8 97 -4
rect 98 -8 102 -4
<< nsubstratencontact >>
rect 21 114 25 118
rect 28 114 32 118
rect 33 114 37 118
rect 38 114 42 118
rect 43 114 47 118
rect 48 114 52 118
rect 53 114 57 118
rect 58 114 62 118
rect 63 114 67 118
rect 68 114 72 118
rect 73 114 77 118
rect 78 114 82 118
rect 85 114 89 118
rect 21 107 25 111
rect 85 107 89 111
rect 21 102 25 106
rect 21 97 25 101
rect 21 92 25 96
rect 21 87 25 91
rect 21 82 25 86
rect 21 77 25 81
rect 21 72 25 76
rect 21 67 25 71
rect 21 62 25 66
rect 21 57 25 61
rect 21 52 25 56
rect 21 47 25 51
rect 21 42 25 46
rect 21 37 25 41
rect 21 32 25 36
rect 21 27 25 31
rect 21 22 25 26
rect 21 17 25 21
rect 85 102 89 106
rect 85 97 89 101
rect 85 92 89 96
rect 85 87 89 91
rect 85 82 89 86
rect 85 77 89 81
rect 85 72 89 76
rect 85 67 89 71
rect 85 62 89 66
rect 85 57 89 61
rect 85 52 89 56
rect 85 47 89 51
rect 85 42 89 46
rect 85 37 89 41
rect 85 32 89 36
rect 85 27 89 31
rect 85 22 89 26
rect 85 17 89 21
rect 21 12 25 16
rect 85 12 89 16
rect 21 5 25 9
rect 28 5 32 9
rect 33 5 37 9
rect 38 5 42 9
rect 43 5 47 9
rect 48 5 52 9
rect 53 5 57 9
rect 58 5 62 9
rect 63 5 67 9
rect 68 5 72 9
rect 73 5 77 9
rect 78 5 82 9
rect 85 5 89 9
<< metal1 >>
rect 12 127 13 131
rect 17 127 18 131
rect 22 127 23 131
rect 27 127 28 131
rect 32 127 33 131
rect 37 127 38 131
rect 42 127 43 131
rect 47 127 48 131
rect 52 127 53 131
rect 57 127 58 131
rect 62 127 63 131
rect 67 127 68 131
rect 72 127 73 131
rect 77 127 78 131
rect 82 127 83 131
rect 87 127 88 131
rect 92 127 93 131
rect 97 127 98 131
rect 8 126 12 127
rect 8 121 12 122
rect 98 126 102 127
rect 98 121 102 122
rect 8 116 12 117
rect 8 111 12 112
rect 8 106 12 107
rect 8 101 12 102
rect 8 96 12 97
rect 8 91 12 92
rect 8 86 12 87
rect 8 81 12 82
rect 8 76 12 77
rect 8 71 12 72
rect 8 66 12 67
rect 8 61 12 62
rect 8 56 12 57
rect 8 51 12 52
rect 8 46 12 47
rect 8 41 12 42
rect 8 36 12 37
rect 8 31 12 32
rect 8 26 12 27
rect 8 21 12 22
rect 8 16 12 17
rect 8 11 12 12
rect 8 6 12 7
rect 25 114 28 118
rect 32 114 33 118
rect 37 114 38 118
rect 42 114 43 118
rect 47 114 48 118
rect 52 114 53 118
rect 57 114 58 118
rect 62 114 63 118
rect 67 114 68 118
rect 72 114 73 118
rect 77 114 78 118
rect 82 114 85 118
rect 21 111 25 114
rect 21 106 25 107
rect 85 111 89 114
rect 85 106 89 107
rect 21 101 25 102
rect 21 96 25 97
rect 21 91 25 92
rect 21 86 25 87
rect 21 81 25 82
rect 21 76 25 77
rect 21 71 25 72
rect 21 66 25 67
rect 21 61 25 62
rect 21 56 25 57
rect 21 51 25 52
rect 21 46 25 47
rect 21 41 25 42
rect 21 36 25 37
rect 21 31 25 32
rect 21 26 25 27
rect 21 21 25 22
rect 32 102 33 106
rect 37 102 38 106
rect 42 102 43 106
rect 47 102 48 106
rect 52 102 53 106
rect 57 102 58 106
rect 62 102 63 106
rect 67 102 68 106
rect 72 102 73 106
rect 32 101 77 102
rect 32 97 33 101
rect 37 97 38 101
rect 42 97 43 101
rect 47 97 48 101
rect 52 97 53 101
rect 57 97 58 101
rect 62 97 63 101
rect 67 97 68 101
rect 72 97 73 101
rect 32 96 77 97
rect 32 92 33 96
rect 37 92 38 96
rect 42 92 43 96
rect 47 92 48 96
rect 52 92 53 96
rect 57 92 58 96
rect 62 92 63 96
rect 67 92 68 96
rect 72 92 73 96
rect 32 91 77 92
rect 32 87 33 91
rect 37 87 38 91
rect 42 87 43 91
rect 47 87 48 91
rect 52 87 53 91
rect 57 87 58 91
rect 62 87 63 91
rect 67 87 68 91
rect 72 87 73 91
rect 32 86 77 87
rect 32 82 33 86
rect 37 82 38 86
rect 42 82 43 86
rect 47 82 48 86
rect 52 82 53 86
rect 57 82 58 86
rect 62 82 63 86
rect 67 82 68 86
rect 72 82 73 86
rect 32 81 77 82
rect 32 77 33 81
rect 37 77 38 81
rect 42 77 43 81
rect 47 77 48 81
rect 52 77 53 81
rect 57 77 58 81
rect 62 77 63 81
rect 67 77 68 81
rect 72 77 73 81
rect 32 76 77 77
rect 32 72 33 76
rect 37 72 38 76
rect 42 72 43 76
rect 47 72 48 76
rect 52 72 53 76
rect 57 72 58 76
rect 62 72 63 76
rect 67 72 68 76
rect 72 72 73 76
rect 32 71 77 72
rect 32 67 33 71
rect 37 67 38 71
rect 42 67 43 71
rect 47 67 48 71
rect 52 67 53 71
rect 57 67 58 71
rect 62 67 63 71
rect 67 67 68 71
rect 72 67 73 71
rect 32 66 77 67
rect 32 62 33 66
rect 37 62 38 66
rect 42 62 43 66
rect 47 62 48 66
rect 52 62 53 66
rect 57 62 58 66
rect 62 62 63 66
rect 67 62 68 66
rect 72 62 73 66
rect 32 61 77 62
rect 32 57 33 61
rect 37 57 38 61
rect 42 57 43 61
rect 47 57 48 61
rect 52 57 53 61
rect 57 57 58 61
rect 62 57 63 61
rect 67 57 68 61
rect 72 57 73 61
rect 32 56 77 57
rect 32 52 33 56
rect 37 52 38 56
rect 42 52 43 56
rect 47 52 48 56
rect 52 52 53 56
rect 57 52 58 56
rect 62 52 63 56
rect 67 52 68 56
rect 72 52 73 56
rect 32 51 77 52
rect 32 47 33 51
rect 37 47 38 51
rect 42 47 43 51
rect 47 47 48 51
rect 52 47 53 51
rect 57 47 58 51
rect 62 47 63 51
rect 67 47 68 51
rect 72 47 73 51
rect 32 46 77 47
rect 32 42 33 46
rect 37 42 38 46
rect 42 42 43 46
rect 47 42 48 46
rect 52 42 53 46
rect 57 42 58 46
rect 62 42 63 46
rect 67 42 68 46
rect 72 42 73 46
rect 32 41 77 42
rect 32 37 33 41
rect 37 37 38 41
rect 42 37 43 41
rect 47 37 48 41
rect 52 37 53 41
rect 57 37 58 41
rect 62 37 63 41
rect 67 37 68 41
rect 72 37 73 41
rect 32 36 77 37
rect 32 32 33 36
rect 37 32 38 36
rect 42 32 43 36
rect 47 32 48 36
rect 52 32 53 36
rect 57 32 58 36
rect 62 32 63 36
rect 67 32 68 36
rect 72 32 73 36
rect 32 31 77 32
rect 32 27 33 31
rect 37 27 38 31
rect 42 27 43 31
rect 47 27 48 31
rect 52 27 53 31
rect 57 27 58 31
rect 62 27 63 31
rect 67 27 68 31
rect 72 27 73 31
rect 32 26 77 27
rect 32 22 33 26
rect 37 22 38 26
rect 42 22 43 26
rect 47 22 48 26
rect 52 22 53 26
rect 57 22 58 26
rect 62 22 63 26
rect 67 22 68 26
rect 72 22 73 26
rect 32 21 77 22
rect 32 17 33 21
rect 37 17 38 21
rect 42 17 43 21
rect 47 17 48 21
rect 52 17 53 21
rect 57 17 58 21
rect 62 17 63 21
rect 67 17 68 21
rect 72 17 73 21
rect 85 101 89 102
rect 85 96 89 97
rect 85 91 89 92
rect 85 86 89 87
rect 85 81 89 82
rect 85 76 89 77
rect 85 71 89 72
rect 85 66 89 67
rect 85 61 89 62
rect 85 56 89 57
rect 85 51 89 52
rect 85 46 89 47
rect 85 41 89 42
rect 85 36 89 37
rect 85 31 89 32
rect 85 26 89 27
rect 85 21 89 22
rect 21 16 25 17
rect 21 9 25 12
rect 85 16 89 17
rect 85 9 89 12
rect 25 5 28 9
rect 32 5 33 9
rect 37 5 38 9
rect 42 5 43 9
rect 47 5 48 9
rect 52 5 53 9
rect 57 5 58 9
rect 62 5 63 9
rect 67 5 68 9
rect 72 5 73 9
rect 77 5 78 9
rect 82 5 85 9
rect 98 116 102 117
rect 98 111 102 112
rect 98 106 102 107
rect 98 101 102 102
rect 98 96 102 97
rect 98 91 102 92
rect 98 86 102 87
rect 98 81 102 82
rect 98 76 102 77
rect 98 71 102 72
rect 98 66 102 67
rect 98 61 102 62
rect 98 56 102 57
rect 98 51 102 52
rect 98 46 102 47
rect 98 41 102 42
rect 98 36 102 37
rect 98 31 102 32
rect 98 26 102 27
rect 98 21 102 22
rect 98 16 102 17
rect 98 11 102 12
rect 98 6 102 7
rect 8 1 12 2
rect 8 -4 12 -3
rect 98 1 102 2
rect 98 -4 102 -3
rect 12 -8 13 -4
rect 17 -8 18 -4
rect 22 -8 23 -4
rect 27 -8 28 -4
rect 32 -8 33 -4
rect 37 -8 38 -4
rect 42 -8 43 -4
rect 47 -8 48 -4
rect 52 -8 53 -4
rect 57 -8 58 -4
rect 62 -8 63 -4
rect 67 -8 68 -4
rect 72 -8 73 -4
rect 77 -8 78 -4
rect 82 -8 83 -4
rect 87 -8 88 -4
rect 92 -8 93 -4
rect 97 -8 98 -4
<< m2contact >>
rect 33 102 37 106
rect 43 102 47 106
rect 53 102 57 106
rect 63 102 67 106
rect 73 102 77 106
rect 38 97 42 101
rect 48 97 52 101
rect 58 97 62 101
rect 68 97 72 101
rect 33 92 37 96
rect 43 92 47 96
rect 53 92 57 96
rect 63 92 67 96
rect 73 92 77 96
rect 38 87 42 91
rect 48 87 52 91
rect 58 87 62 91
rect 68 87 72 91
rect 33 82 37 86
rect 43 82 47 86
rect 53 82 57 86
rect 63 82 67 86
rect 73 82 77 86
rect 38 77 42 81
rect 48 77 52 81
rect 58 77 62 81
rect 68 77 72 81
rect 33 72 37 76
rect 43 72 47 76
rect 53 72 57 76
rect 63 72 67 76
rect 73 72 77 76
rect 38 67 42 71
rect 48 67 52 71
rect 58 67 62 71
rect 68 67 72 71
rect 33 62 37 66
rect 43 62 47 66
rect 53 62 57 66
rect 63 62 67 66
rect 73 62 77 66
rect 38 57 42 61
rect 48 57 52 61
rect 58 57 62 61
rect 68 57 72 61
rect 33 52 37 56
rect 43 52 47 56
rect 53 52 57 56
rect 63 52 67 56
rect 73 52 77 56
rect 38 47 42 51
rect 48 47 52 51
rect 58 47 62 51
rect 68 47 72 51
rect 33 42 37 46
rect 43 42 47 46
rect 53 42 57 46
rect 63 42 67 46
rect 73 42 77 46
rect 38 37 42 41
rect 48 37 52 41
rect 58 37 62 41
rect 68 37 72 41
rect 33 32 37 36
rect 43 32 47 36
rect 53 32 57 36
rect 63 32 67 36
rect 73 32 77 36
rect 38 27 42 31
rect 48 27 52 31
rect 58 27 62 31
rect 68 27 72 31
rect 33 22 37 26
rect 43 22 47 26
rect 53 22 57 26
rect 63 22 67 26
rect 73 22 77 26
rect 38 17 42 21
rect 48 17 52 21
rect 58 17 62 21
rect 68 17 72 21
<< metal2 >>
rect 37 102 43 106
rect 47 102 53 106
rect 57 102 63 106
rect 67 102 73 106
rect 33 101 77 102
rect 33 97 38 101
rect 42 97 48 101
rect 52 97 58 101
rect 62 97 68 101
rect 72 97 77 101
rect 33 96 77 97
rect 37 92 43 96
rect 47 92 53 96
rect 57 92 63 96
rect 67 92 73 96
rect 33 91 77 92
rect 33 87 38 91
rect 42 87 48 91
rect 52 87 58 91
rect 62 87 68 91
rect 72 87 77 91
rect 33 86 77 87
rect 37 82 43 86
rect 47 82 53 86
rect 57 82 63 86
rect 67 82 73 86
rect 33 81 77 82
rect 33 77 38 81
rect 42 77 48 81
rect 52 77 58 81
rect 62 77 68 81
rect 72 77 77 81
rect 33 76 77 77
rect 37 72 43 76
rect 47 72 53 76
rect 57 72 63 76
rect 67 72 73 76
rect 33 71 77 72
rect 33 67 38 71
rect 42 67 48 71
rect 52 67 58 71
rect 62 67 68 71
rect 72 67 77 71
rect 33 66 77 67
rect 37 62 43 66
rect 47 62 53 66
rect 57 62 63 66
rect 67 62 73 66
rect 33 61 77 62
rect 33 57 38 61
rect 42 57 48 61
rect 52 57 58 61
rect 62 57 68 61
rect 72 57 77 61
rect 33 56 77 57
rect 37 52 43 56
rect 47 52 53 56
rect 57 52 63 56
rect 67 52 73 56
rect 33 51 77 52
rect 33 47 38 51
rect 42 47 48 51
rect 52 47 58 51
rect 62 47 68 51
rect 72 47 77 51
rect 33 46 77 47
rect 37 42 43 46
rect 47 42 53 46
rect 57 42 63 46
rect 67 42 73 46
rect 33 41 77 42
rect 33 37 38 41
rect 42 37 48 41
rect 52 37 58 41
rect 62 37 68 41
rect 72 37 77 41
rect 33 36 77 37
rect 37 32 43 36
rect 47 32 53 36
rect 57 32 63 36
rect 67 32 73 36
rect 33 31 77 32
rect 33 27 38 31
rect 42 27 48 31
rect 52 27 58 31
rect 62 27 68 31
rect 72 27 77 31
rect 33 26 77 27
rect 37 22 43 26
rect 47 22 53 26
rect 57 22 63 26
rect 67 22 73 26
rect 33 21 77 22
rect 33 17 38 21
rect 42 17 48 21
rect 52 17 58 21
rect 62 17 68 21
rect 72 17 77 21
<< end >>
