magic
tech scmos
timestamp 1012172318
<< ntransistor >>
rect 193 313 252 315
rect 193 305 252 307
rect 193 297 252 299
rect 193 289 252 291
rect 193 272 252 274
rect 193 264 252 266
rect 193 256 252 258
rect 193 248 252 250
rect 193 229 252 231
rect 193 221 252 223
rect 193 213 252 215
rect 193 205 252 207
rect 193 190 233 192
rect 193 182 233 184
rect 193 174 233 176
rect 193 166 233 168
rect 193 158 233 160
rect 193 150 233 152
<< ptransistor >>
rect 75 313 163 315
rect 75 305 163 307
rect 75 297 163 299
rect 75 289 163 291
rect 75 272 163 274
rect 75 264 163 266
rect 75 256 163 258
rect 75 248 163 250
rect 75 229 163 231
rect 75 221 163 223
rect 75 213 163 215
rect 75 205 163 207
rect 107 190 163 192
rect 107 182 163 184
rect 107 174 163 176
rect 107 166 163 168
rect 107 158 163 160
rect 107 150 163 152
<< ndiffusion >>
rect 193 320 252 321
rect 200 316 204 320
rect 193 315 252 316
rect 193 312 252 313
rect 193 307 252 308
rect 193 304 252 305
rect 193 300 204 304
rect 193 299 252 300
rect 193 296 252 297
rect 193 291 252 292
rect 193 284 252 289
rect 193 279 252 280
rect 200 275 204 279
rect 193 274 252 275
rect 193 271 252 272
rect 193 266 252 267
rect 193 263 252 264
rect 193 259 204 263
rect 193 258 252 259
rect 193 255 252 256
rect 193 250 252 251
rect 193 241 252 248
rect 193 236 252 237
rect 200 232 204 236
rect 193 231 252 232
rect 193 228 252 229
rect 193 223 252 224
rect 193 220 252 221
rect 200 216 204 220
rect 193 215 252 216
rect 193 212 252 213
rect 193 207 252 208
rect 193 202 252 205
rect 193 197 233 198
rect 200 193 204 197
rect 193 192 233 193
rect 193 189 233 190
rect 193 184 233 185
rect 193 181 233 182
rect 200 177 204 181
rect 193 176 233 177
rect 193 173 233 174
rect 193 168 233 169
rect 193 165 233 166
rect 200 161 204 165
rect 193 160 233 161
rect 193 157 233 158
rect 193 152 233 153
rect 193 149 233 150
rect 200 145 204 149
<< pdiffusion >>
rect 75 320 163 321
rect 142 316 146 320
rect 75 315 163 316
rect 75 312 163 313
rect 75 307 163 308
rect 75 304 163 305
rect 142 300 146 304
rect 154 300 163 304
rect 75 299 163 300
rect 75 296 163 297
rect 75 291 163 292
rect 75 284 163 289
rect 75 279 163 280
rect 142 275 146 279
rect 75 274 163 275
rect 75 271 163 272
rect 75 266 163 267
rect 75 263 163 264
rect 142 259 146 263
rect 154 259 163 263
rect 75 258 163 259
rect 75 255 163 256
rect 75 250 163 251
rect 75 245 163 248
rect 75 236 163 237
rect 142 232 146 236
rect 75 231 163 232
rect 75 228 163 229
rect 75 223 163 224
rect 75 220 163 221
rect 142 216 146 220
rect 154 216 163 220
rect 75 215 163 216
rect 75 212 163 213
rect 75 207 163 208
rect 75 202 163 205
rect 107 197 163 198
rect 142 193 146 197
rect 107 192 163 193
rect 107 189 163 190
rect 107 184 163 185
rect 107 181 163 182
rect 142 177 146 181
rect 107 176 163 177
rect 107 173 163 174
rect 107 168 163 169
rect 107 165 163 166
rect 142 161 146 165
rect 107 160 163 161
rect 107 157 163 158
rect 107 152 163 153
rect 107 149 163 150
rect 142 145 146 149
<< ndcontact >>
rect 193 316 200 320
rect 204 316 252 320
rect 193 308 252 312
rect 204 300 252 304
rect 193 292 252 296
rect 193 275 200 279
rect 204 275 252 279
rect 193 267 252 271
rect 204 259 252 263
rect 193 251 252 255
rect 193 232 200 236
rect 204 232 252 236
rect 193 224 252 228
rect 193 216 200 220
rect 204 216 252 220
rect 193 208 252 212
rect 193 193 200 197
rect 204 193 233 197
rect 193 185 233 189
rect 193 177 200 181
rect 204 177 233 181
rect 193 169 233 173
rect 193 161 200 165
rect 204 161 233 165
rect 193 153 233 157
rect 193 145 200 149
rect 204 145 233 149
<< pdcontact >>
rect 75 316 142 320
rect 146 316 163 320
rect 75 308 163 312
rect 75 300 142 304
rect 146 300 154 304
rect 75 292 163 296
rect 75 275 142 279
rect 146 275 163 279
rect 75 267 163 271
rect 75 259 142 263
rect 146 259 154 263
rect 75 251 163 255
rect 75 232 142 236
rect 146 232 163 236
rect 75 224 163 228
rect 75 216 142 220
rect 146 216 154 220
rect 75 208 163 212
rect 107 193 142 197
rect 146 193 163 197
rect 107 185 163 189
rect 107 177 142 181
rect 146 177 163 181
rect 107 169 163 173
rect 107 161 142 165
rect 146 161 163 165
rect 107 153 163 157
rect 107 145 142 149
rect 146 145 163 149
<< psubstratepcontact >>
rect 193 321 252 325
rect 193 280 252 284
rect 193 237 252 241
rect 193 198 233 202
<< nsubstratencontact >>
rect 75 321 163 325
rect 75 280 163 284
rect 75 237 163 241
rect 107 198 163 202
<< polysilicon >>
rect 72 313 75 315
rect 163 313 193 315
rect 252 313 255 315
rect 72 307 74 313
rect 166 307 192 313
rect 253 307 255 313
rect 72 305 75 307
rect 163 305 193 307
rect 252 305 255 307
rect 72 299 74 305
rect 166 299 192 305
rect 72 297 75 299
rect 163 297 193 299
rect 252 297 255 299
rect 72 291 74 297
rect 166 291 192 297
rect 253 291 255 297
rect 72 289 75 291
rect 163 289 193 291
rect 252 289 255 291
rect 168 288 192 289
rect 168 282 172 288
rect 181 282 192 288
rect 168 274 192 282
rect 72 272 75 274
rect 163 272 193 274
rect 252 272 255 274
rect 72 266 74 272
rect 166 266 192 272
rect 253 266 255 272
rect 72 264 75 266
rect 163 264 193 266
rect 252 264 255 266
rect 72 258 74 264
rect 166 258 192 264
rect 72 256 75 258
rect 163 256 193 258
rect 252 256 255 258
rect 72 250 74 256
rect 166 253 192 256
rect 166 250 170 253
rect 72 248 75 250
rect 163 249 170 250
rect 183 250 192 253
rect 253 250 255 256
rect 183 249 193 250
rect 163 248 193 249
rect 252 248 255 250
rect 72 229 75 231
rect 163 229 166 231
rect 72 223 74 229
rect 164 223 166 229
rect 72 221 75 223
rect 163 221 166 223
rect 72 215 74 221
rect 164 215 166 221
rect 72 213 75 215
rect 163 213 166 215
rect 72 207 74 213
rect 164 212 166 213
rect 190 229 193 231
rect 252 229 255 231
rect 190 223 192 229
rect 253 223 255 229
rect 190 221 193 223
rect 252 221 255 223
rect 190 215 192 221
rect 190 213 193 215
rect 252 213 255 215
rect 190 212 192 213
rect 164 210 192 212
rect 164 207 168 210
rect 72 205 75 207
rect 163 206 168 207
rect 181 207 192 210
rect 253 207 255 213
rect 181 206 193 207
rect 163 205 193 206
rect 252 205 255 207
rect 104 190 107 192
rect 163 190 166 192
rect 104 184 106 190
rect 164 184 166 190
rect 104 182 107 184
rect 163 182 166 184
rect 104 176 106 182
rect 164 176 166 182
rect 104 174 107 176
rect 163 174 166 176
rect 104 168 106 174
rect 164 170 166 174
rect 190 190 193 192
rect 233 190 236 192
rect 190 184 192 190
rect 234 184 236 190
rect 190 182 193 184
rect 233 182 236 184
rect 190 176 192 182
rect 234 176 236 182
rect 190 174 193 176
rect 233 174 236 176
rect 190 170 192 174
rect 164 168 192 170
rect 234 168 236 174
rect 104 166 107 168
rect 163 166 177 168
rect 183 166 193 168
rect 233 166 236 168
rect 105 158 107 160
rect 163 158 193 160
rect 233 158 235 160
rect 170 152 172 158
rect 105 150 107 152
rect 163 150 193 152
rect 233 150 235 152
rect 172 147 178 150
<< polycontact >>
rect 172 282 181 288
rect 170 249 183 253
rect 168 206 181 210
rect 177 164 183 168
rect 172 143 178 147
<< metal1 >>
rect 114 357 230 366
rect 124 345 220 357
rect 48 321 75 325
rect 48 320 163 321
rect 48 316 75 320
rect 48 304 72 316
rect 170 312 188 345
rect 252 321 298 325
rect 193 320 298 321
rect 252 316 298 320
rect 163 308 193 312
rect 48 300 75 304
rect 48 284 72 300
rect 157 296 193 308
rect 257 304 298 316
rect 252 300 298 304
rect 163 292 193 296
rect 48 280 75 284
rect 48 279 163 280
rect 48 275 75 279
rect 48 263 72 275
rect 184 271 190 292
rect 257 284 298 300
rect 252 280 298 284
rect 193 279 298 280
rect 252 275 298 279
rect 163 267 193 271
rect 48 259 75 263
rect 157 262 192 267
rect 257 263 298 275
rect 48 241 72 259
rect 157 255 163 262
rect 188 255 192 262
rect 252 259 298 263
rect 170 253 183 254
rect 188 251 193 255
rect 48 237 75 241
rect 48 236 163 237
rect 48 232 75 236
rect 170 238 183 249
rect 257 241 298 259
rect 48 220 72 232
rect 170 230 172 238
rect 181 230 183 238
rect 252 237 298 241
rect 193 236 298 237
rect 252 232 298 236
rect 170 228 183 230
rect 163 224 193 228
rect 48 216 75 220
rect 157 219 190 224
rect 255 220 298 232
rect 48 197 72 216
rect 157 212 163 219
rect 186 212 190 219
rect 252 216 298 220
rect 168 210 181 211
rect 186 208 193 212
rect 107 197 163 198
rect 48 193 107 197
rect 48 181 104 193
rect 168 189 181 206
rect 193 197 233 198
rect 255 197 298 216
rect 233 193 298 197
rect 163 185 193 189
rect 48 177 107 181
rect 48 166 104 177
rect 167 176 190 185
rect 242 181 298 193
rect 233 177 298 181
rect 167 173 174 176
rect 163 169 174 173
rect 186 173 190 176
rect 186 169 193 173
rect 36 165 104 166
rect 36 164 107 165
rect 36 160 37 164
rect 41 160 42 164
rect 46 161 107 164
rect 242 165 298 177
rect 46 160 104 161
rect 36 159 104 160
rect 36 155 37 159
rect 41 155 42 159
rect 46 155 104 159
rect 177 157 181 164
rect 233 161 298 165
rect 36 154 104 155
rect 36 150 37 154
rect 41 150 42 154
rect 46 150 104 154
rect 163 153 193 157
rect 36 149 104 150
rect 242 149 298 161
rect 36 145 37 149
rect 41 145 42 149
rect 46 145 107 149
rect 36 144 104 145
rect 36 140 37 144
rect 41 140 42 144
rect 46 140 104 144
rect 233 145 298 149
rect 36 139 104 140
rect 36 135 37 139
rect 41 135 42 139
rect 46 135 104 139
rect 36 134 104 135
rect 36 130 37 134
rect 41 130 42 134
rect 46 130 104 134
rect 36 129 104 130
rect 36 125 37 129
rect 41 125 42 129
rect 46 125 104 129
rect 36 124 104 125
rect 36 120 37 124
rect 41 120 42 124
rect 46 120 104 124
rect 36 119 104 120
rect 36 115 37 119
rect 41 115 42 119
rect 46 115 104 119
rect 36 114 104 115
rect 36 110 37 114
rect 41 110 42 114
rect 46 110 104 114
rect 36 109 104 110
rect 36 105 37 109
rect 41 105 42 109
rect 46 105 104 109
rect 36 104 104 105
rect 36 100 37 104
rect 41 100 42 104
rect 46 100 104 104
rect 36 98 104 100
rect 168 -26 181 143
rect 242 86 298 145
rect 246 82 247 86
rect 251 82 252 86
rect 256 82 257 86
rect 261 82 262 86
rect 266 82 267 86
rect 271 82 272 86
rect 276 82 277 86
rect 281 82 282 86
rect 286 82 287 86
rect 291 82 292 86
rect 296 82 298 86
rect 242 81 298 82
rect 246 77 247 81
rect 251 77 252 81
rect 256 77 257 81
rect 261 77 262 81
rect 266 77 267 81
rect 271 77 272 81
rect 276 77 277 81
rect 281 77 282 81
rect 286 77 287 81
rect 291 77 292 81
rect 296 77 298 81
rect 242 76 298 77
<< m2contact >>
rect 142 316 146 320
rect 200 316 204 320
rect 142 300 146 304
rect 200 300 204 304
rect 142 275 146 279
rect 172 274 181 282
rect 200 275 204 279
rect 142 259 146 263
rect 200 259 204 263
rect 142 232 146 236
rect 172 230 181 238
rect 200 232 204 236
rect 142 216 146 220
rect 200 216 204 220
rect 142 193 146 197
rect 200 193 204 197
rect 142 177 146 181
rect 200 177 204 181
rect 37 160 41 164
rect 42 160 46 164
rect 142 161 146 165
rect 37 155 41 159
rect 42 155 46 159
rect 200 161 204 165
rect 37 150 41 154
rect 42 150 46 154
rect 37 145 41 149
rect 42 145 46 149
rect 142 145 146 149
rect 37 140 41 144
rect 42 140 46 144
rect 200 145 204 149
rect 37 135 41 139
rect 42 135 46 139
rect 37 130 41 134
rect 42 130 46 134
rect 37 125 41 129
rect 42 125 46 129
rect 37 120 41 124
rect 42 120 46 124
rect 37 115 41 119
rect 42 115 46 119
rect 37 110 41 114
rect 42 110 46 114
rect 37 105 41 109
rect 42 105 46 109
rect 37 100 41 104
rect 42 100 46 104
rect 242 82 246 86
rect 247 82 251 86
rect 252 82 256 86
rect 257 82 261 86
rect 262 82 266 86
rect 267 82 271 86
rect 272 82 276 86
rect 277 82 281 86
rect 282 82 286 86
rect 287 82 291 86
rect 292 82 296 86
rect 242 77 246 81
rect 247 77 251 81
rect 252 77 256 81
rect 257 77 261 81
rect 262 77 266 81
rect 267 77 271 81
rect 272 77 276 81
rect 277 77 281 81
rect 282 77 286 81
rect 287 77 291 81
rect 292 77 296 81
<< metal2 >>
rect 142 304 146 316
rect 142 279 146 300
rect 200 304 204 316
rect 142 263 146 275
rect 142 236 146 259
rect 142 220 146 232
rect 170 282 183 288
rect 170 274 172 282
rect 181 274 183 282
rect 170 238 183 274
rect 170 230 172 238
rect 181 230 183 238
rect 170 228 183 230
rect 200 279 204 300
rect 200 263 204 275
rect 200 236 204 259
rect 142 197 146 216
rect 142 181 146 193
rect 25 164 46 166
rect 25 160 27 164
rect 31 160 32 164
rect 36 160 37 164
rect 41 160 42 164
rect 25 159 46 160
rect 25 155 27 159
rect 31 155 32 159
rect 36 155 37 159
rect 41 155 42 159
rect 25 154 46 155
rect 25 150 27 154
rect 31 150 32 154
rect 36 150 37 154
rect 41 150 42 154
rect 25 149 46 150
rect 25 145 27 149
rect 31 145 32 149
rect 36 145 37 149
rect 41 145 42 149
rect 142 165 146 177
rect 142 149 146 161
rect 200 220 204 232
rect 200 197 204 216
rect 200 181 204 193
rect 200 165 204 177
rect 200 149 204 161
rect 25 144 46 145
rect 25 140 27 144
rect 31 140 32 144
rect 36 140 37 144
rect 41 140 42 144
rect 25 139 46 140
rect 25 135 27 139
rect 31 135 32 139
rect 36 135 37 139
rect 41 135 42 139
rect 25 134 46 135
rect 25 130 27 134
rect 31 130 32 134
rect 36 130 37 134
rect 41 130 42 134
rect 25 129 46 130
rect 25 125 27 129
rect 31 125 32 129
rect 36 125 37 129
rect 41 125 42 129
rect 25 124 46 125
rect 25 120 27 124
rect 31 120 32 124
rect 36 120 37 124
rect 41 120 42 124
rect 25 119 46 120
rect 25 115 27 119
rect 31 115 32 119
rect 36 115 37 119
rect 41 115 42 119
rect 25 114 46 115
rect 25 110 27 114
rect 31 110 32 114
rect 36 110 37 114
rect 41 110 42 114
rect 25 109 46 110
rect 25 105 27 109
rect 31 105 32 109
rect 36 105 37 109
rect 41 105 42 109
rect 25 104 46 105
rect 25 100 27 104
rect 31 100 32 104
rect 36 100 37 104
rect 41 100 42 104
rect 25 98 46 100
rect 246 82 247 86
rect 251 82 252 86
rect 256 82 257 86
rect 261 82 262 86
rect 266 82 267 86
rect 271 82 272 86
rect 276 82 277 86
rect 281 82 282 86
rect 286 82 287 86
rect 291 82 292 86
rect 296 82 298 86
rect 242 81 298 82
rect 246 77 247 81
rect 251 77 252 81
rect 256 77 257 81
rect 261 77 262 81
rect 266 77 267 81
rect 271 77 272 81
rect 276 77 277 81
rect 281 77 282 81
rect 286 77 287 81
rect 291 77 292 81
rect 296 77 298 81
rect 242 76 298 77
rect 246 72 247 76
rect 251 72 252 76
rect 256 72 257 76
rect 261 72 262 76
rect 266 72 267 76
rect 271 72 272 76
rect 276 72 277 76
rect 281 72 282 76
rect 286 72 287 76
rect 291 72 292 76
rect 296 72 298 76
rect 242 71 298 72
rect 246 67 247 71
rect 251 67 252 71
rect 256 67 257 71
rect 261 67 262 71
rect 266 67 267 71
rect 271 67 272 71
rect 276 67 277 71
rect 281 67 282 71
rect 286 67 287 71
rect 291 67 292 71
rect 296 67 298 71
rect 242 65 298 67
<< m3contact >>
rect 27 160 31 164
rect 32 160 36 164
rect 27 155 31 159
rect 32 155 36 159
rect 27 150 31 154
rect 32 150 36 154
rect 27 145 31 149
rect 32 145 36 149
rect 27 140 31 144
rect 32 140 36 144
rect 27 135 31 139
rect 32 135 36 139
rect 27 130 31 134
rect 32 130 36 134
rect 27 125 31 129
rect 32 125 36 129
rect 27 120 31 124
rect 32 120 36 124
rect 27 115 31 119
rect 32 115 36 119
rect 27 110 31 114
rect 32 110 36 114
rect 27 105 31 109
rect 32 105 36 109
rect 27 100 31 104
rect 32 100 36 104
rect 242 72 246 76
rect 247 72 251 76
rect 252 72 256 76
rect 257 72 261 76
rect 262 72 266 76
rect 267 72 271 76
rect 272 72 276 76
rect 277 72 281 76
rect 282 72 286 76
rect 287 72 291 76
rect 292 72 296 76
rect 242 67 246 71
rect 247 67 251 71
rect 252 67 256 71
rect 257 67 261 71
rect 262 67 266 71
rect 267 67 271 71
rect 272 67 276 71
rect 277 67 281 71
rect 282 67 286 71
rect 287 67 291 71
rect 292 67 296 71
<< metal3 >>
rect 25 164 37 166
rect 25 160 27 164
rect 31 160 32 164
rect 36 160 37 164
rect 25 159 37 160
rect 25 155 27 159
rect 31 155 32 159
rect 36 155 37 159
rect 25 154 37 155
rect 25 150 27 154
rect 31 150 32 154
rect 36 150 37 154
rect 25 149 37 150
rect 25 145 27 149
rect 31 145 32 149
rect 36 145 37 149
rect 25 144 37 145
rect 25 140 27 144
rect 31 140 32 144
rect 36 140 37 144
rect 25 139 37 140
rect 25 135 27 139
rect 31 135 32 139
rect 36 135 37 139
rect 25 134 37 135
rect 25 130 27 134
rect 31 130 32 134
rect 36 130 37 134
rect 25 129 37 130
rect 25 125 27 129
rect 31 125 32 129
rect 36 125 37 129
rect 25 124 37 125
rect 25 120 27 124
rect 31 120 32 124
rect 36 120 37 124
rect 25 119 37 120
rect 25 115 27 119
rect 31 115 32 119
rect 36 115 37 119
rect 25 114 37 115
rect 25 110 27 114
rect 31 110 32 114
rect 36 110 37 114
rect 25 109 37 110
rect 25 105 27 109
rect 31 105 32 109
rect 36 105 37 109
rect 25 104 37 105
rect 25 100 27 104
rect 31 100 32 104
rect 36 100 37 104
rect 25 97 37 100
rect 241 76 298 78
rect 241 72 242 76
rect 246 72 247 76
rect 251 72 252 76
rect 256 72 257 76
rect 261 72 262 76
rect 266 72 267 76
rect 271 72 272 76
rect 276 72 277 76
rect 281 72 282 76
rect 286 72 287 76
rect 291 72 292 76
rect 296 72 298 76
rect 241 71 298 72
rect 241 67 242 71
rect 246 67 247 71
rect 251 67 252 71
rect 256 67 257 71
rect 261 67 262 71
rect 266 67 267 71
rect 271 67 272 71
rect 276 67 277 71
rect 281 67 282 71
rect 286 67 287 71
rect 291 67 292 71
rect 296 67 298 71
rect 241 65 298 67
use barepad b
timestamp 1006127261
transform 1 0 26 0 1 -357
box 16 702 276 1014
use barering br
timestamp 1006127261
transform 1 0 15 0 1 -3
box 2 -23 311 176
<< labels >>
rlabel metal3 32 103 32 103 1 Vdd!
rlabel metal1 174 12 174 12 1 out
rlabel polycontact 180 166 180 166 1 _out
rlabel metal1 172 352 172 352 1 RawOut
<< end >>
