magic
tech scmos
timestamp 1512385298
<< metal1 >>
rect -9 1974 -5 4676
rect -2 1974 2 4676
rect 5 1974 9 4676
rect 12 1974 16 4676
rect 19 1974 23 4676
rect 26 1974 30 4676
rect 33 1974 37 4676
rect 40 1974 44 4676
rect 47 1974 51 4676
rect 54 1974 58 4676
<< end >>
