magic
tech scmos
timestamp 1509371954
<< ntransistor >>
rect 144 -152 184 -150
rect 144 -160 184 -158
rect 144 -168 184 -166
rect 144 -176 184 -174
rect 144 -184 184 -182
rect 144 -192 184 -190
<< ptransistor >>
rect 58 -152 114 -150
rect 58 -160 114 -158
rect 58 -168 114 -166
rect 58 -176 114 -174
rect 58 -184 114 -182
rect 58 -192 114 -190
<< ndiffusion >>
rect 151 -149 155 -145
rect 144 -150 184 -149
rect 144 -153 184 -152
rect 144 -158 184 -157
rect 144 -161 184 -160
rect 151 -165 155 -161
rect 144 -166 184 -165
rect 144 -169 184 -168
rect 144 -174 184 -173
rect 144 -177 184 -176
rect 151 -181 155 -177
rect 144 -182 184 -181
rect 144 -185 184 -184
rect 144 -190 184 -189
rect 144 -193 184 -192
rect 151 -197 155 -193
<< pdiffusion >>
rect 93 -149 97 -145
rect 58 -150 114 -149
rect 58 -153 114 -152
rect 58 -158 114 -157
rect 58 -161 114 -160
rect 93 -165 97 -161
rect 58 -166 114 -165
rect 58 -169 114 -168
rect 58 -174 114 -173
rect 58 -177 114 -176
rect 93 -181 97 -177
rect 58 -182 114 -181
rect 58 -185 114 -184
rect 58 -190 114 -189
rect 58 -193 114 -192
rect 93 -197 97 -193
<< ndcontact >>
rect 144 -149 151 -145
rect 155 -149 184 -145
rect 144 -157 184 -153
rect 144 -165 151 -161
rect 155 -165 184 -161
rect 144 -173 184 -169
rect 144 -181 151 -177
rect 155 -181 184 -177
rect 144 -189 184 -185
rect 144 -197 151 -193
rect 155 -197 184 -193
<< pdcontact >>
rect 58 -149 93 -145
rect 97 -149 114 -145
rect 58 -157 114 -153
rect 58 -165 93 -161
rect 97 -165 114 -161
rect 58 -173 114 -169
rect 58 -181 93 -177
rect 97 -181 114 -177
rect 58 -189 114 -185
rect 58 -197 93 -193
rect 97 -197 114 -193
<< polysilicon >>
rect 112 -93 133 -24
rect 118 -150 127 -149
rect 56 -152 58 -150
rect 114 -152 144 -150
rect 184 -152 186 -150
rect 121 -158 123 -152
rect 56 -160 58 -158
rect 114 -160 144 -158
rect 184 -160 186 -158
rect 55 -168 58 -166
rect 114 -168 128 -166
rect 134 -168 144 -166
rect 184 -168 187 -166
rect 55 -174 57 -168
rect 115 -170 143 -168
rect 115 -174 117 -170
rect 55 -176 58 -174
rect 114 -176 117 -174
rect 55 -182 57 -176
rect 115 -182 117 -176
rect 55 -184 58 -182
rect 114 -184 117 -182
rect 55 -190 57 -184
rect 115 -190 117 -184
rect 55 -192 58 -190
rect 114 -192 117 -190
rect 141 -174 143 -170
rect 185 -174 187 -168
rect 141 -176 144 -174
rect 184 -176 187 -174
rect 141 -182 143 -176
rect 185 -182 187 -176
rect 141 -184 144 -182
rect 184 -184 187 -182
rect 141 -190 143 -184
rect 185 -190 187 -184
rect 141 -192 144 -190
rect 184 -192 187 -190
<< polycontact >>
rect 112 -24 133 -15
rect 112 -102 133 -93
rect 118 -149 127 -145
rect 128 -168 134 -164
<< metal1 >>
rect 65 25 181 26
rect 65 21 78 25
rect 82 21 85 25
rect 89 21 92 25
rect 96 21 99 25
rect 103 21 106 25
rect 110 21 113 25
rect 117 21 120 25
rect 124 21 127 25
rect 131 21 134 25
rect 138 21 141 25
rect 145 21 148 25
rect 152 21 155 25
rect 159 21 162 25
rect 166 21 181 25
rect 65 20 181 21
rect 65 17 78 20
rect 75 16 78 17
rect 82 16 85 20
rect 89 16 92 20
rect 96 16 99 20
rect 103 16 106 20
rect 110 16 113 20
rect 117 16 120 20
rect 124 16 127 20
rect 131 16 134 20
rect 138 16 141 20
rect 145 16 148 20
rect 152 16 155 20
rect 159 16 162 20
rect 166 17 181 20
rect 166 16 171 17
rect 75 15 171 16
rect 75 11 78 15
rect 82 11 85 15
rect 89 11 92 15
rect 96 11 99 15
rect 103 11 106 15
rect 110 11 113 15
rect 117 11 120 15
rect 124 11 127 15
rect 131 11 134 15
rect 138 11 141 15
rect 145 11 148 15
rect 152 11 155 15
rect 159 11 162 15
rect 166 11 171 15
rect 75 10 171 11
rect 75 6 78 10
rect 82 6 85 10
rect 89 6 92 10
rect 96 6 99 10
rect 103 6 106 10
rect 110 6 113 10
rect 117 6 120 10
rect 124 6 127 10
rect 131 6 134 10
rect 138 6 141 10
rect 145 6 148 10
rect 152 6 155 10
rect 159 6 162 10
rect 166 6 171 10
rect 75 5 171 6
rect 112 -15 133 5
rect 13 -128 16 -124
rect 20 -128 21 -124
rect 25 -128 26 -124
rect 30 -128 31 -124
rect 35 -128 36 -124
rect 40 -128 41 -124
rect 45 -128 46 -124
rect 50 -128 51 -124
rect 55 -128 56 -124
rect 60 -128 61 -124
rect 65 -128 66 -124
rect 70 -128 73 -124
rect 112 -130 133 -102
rect 173 -128 176 -124
rect 180 -128 181 -124
rect 185 -128 186 -124
rect 190 -128 191 -124
rect 195 -128 196 -124
rect 200 -128 201 -124
rect 205 -128 206 -124
rect 210 -128 211 -124
rect 215 -128 216 -124
rect 220 -128 221 -124
rect 225 -128 226 -124
rect 230 -128 233 -124
rect 114 -132 131 -130
rect 116 -134 129 -132
rect -1 -145 55 -137
rect 118 -145 127 -134
rect 193 -145 249 -137
rect -1 -149 58 -145
rect 184 -149 249 -145
rect -1 -161 55 -149
rect 114 -157 144 -153
rect -1 -165 58 -161
rect 128 -164 132 -157
rect 193 -161 249 -149
rect -1 -174 55 -165
rect 184 -165 249 -161
rect 114 -173 125 -169
rect -13 -176 55 -174
rect -13 -180 -12 -176
rect -8 -180 -7 -176
rect -3 -177 55 -176
rect 118 -176 125 -173
rect 137 -173 144 -169
rect 137 -176 141 -173
rect -3 -180 58 -177
rect -13 -181 58 -180
rect -13 -185 -12 -181
rect -8 -185 -7 -181
rect -3 -185 55 -181
rect 118 -185 141 -176
rect 193 -177 249 -165
rect 184 -181 249 -177
rect -13 -186 55 -185
rect -13 -190 -12 -186
rect -8 -190 -7 -186
rect -3 -190 55 -186
rect 114 -189 144 -185
rect -13 -191 55 -190
rect -13 -195 -12 -191
rect -8 -195 -7 -191
rect -3 -193 55 -191
rect -3 -195 58 -193
rect -13 -196 58 -195
rect -13 -200 -12 -196
rect -8 -200 -7 -196
rect -3 -197 58 -196
rect -3 -200 55 -197
rect -13 -201 55 -200
rect -13 -205 -12 -201
rect -8 -205 -7 -201
rect -3 -205 55 -201
rect -13 -206 55 -205
rect -13 -210 -12 -206
rect -8 -210 -7 -206
rect -3 -210 55 -206
rect -13 -211 55 -210
rect -13 -215 -12 -211
rect -8 -215 -7 -211
rect -3 -215 55 -211
rect -13 -216 55 -215
rect -13 -220 -12 -216
rect -8 -220 -7 -216
rect -3 -220 55 -216
rect -13 -221 55 -220
rect -13 -225 -12 -221
rect -8 -225 -7 -221
rect -3 -225 55 -221
rect -13 -226 55 -225
rect -13 -230 -12 -226
rect -8 -230 -7 -226
rect -3 -230 55 -226
rect -13 -231 55 -230
rect -13 -235 -12 -231
rect -8 -235 -7 -231
rect -3 -235 55 -231
rect -13 -236 55 -235
rect -13 -240 -12 -236
rect -8 -240 -7 -236
rect -3 -240 55 -236
rect -13 -242 55 -240
rect 119 -366 132 -189
rect 193 -193 249 -181
rect 184 -197 249 -193
rect 193 -254 249 -197
rect 197 -258 198 -254
rect 202 -258 203 -254
rect 207 -258 208 -254
rect 212 -258 213 -254
rect 217 -258 218 -254
rect 222 -258 223 -254
rect 227 -258 228 -254
rect 232 -258 233 -254
rect 237 -258 238 -254
rect 242 -258 243 -254
rect 247 -258 249 -254
rect 193 -259 249 -258
rect 197 -263 198 -259
rect 202 -263 203 -259
rect 207 -263 208 -259
rect 212 -263 213 -259
rect 217 -263 218 -259
rect 222 -263 223 -259
rect 227 -263 228 -259
rect 232 -263 233 -259
rect 237 -263 238 -259
rect 242 -263 243 -259
rect 247 -263 249 -259
rect 193 -264 249 -263
<< m2contact >>
rect 78 21 82 25
rect 85 21 89 25
rect 92 21 96 25
rect 99 21 103 25
rect 106 21 110 25
rect 113 21 117 25
rect 120 21 124 25
rect 127 21 131 25
rect 134 21 138 25
rect 141 21 145 25
rect 148 21 152 25
rect 155 21 159 25
rect 162 21 166 25
rect 78 16 82 20
rect 85 16 89 20
rect 92 16 96 20
rect 99 16 103 20
rect 106 16 110 20
rect 113 16 117 20
rect 120 16 124 20
rect 127 16 131 20
rect 134 16 138 20
rect 141 16 145 20
rect 148 16 152 20
rect 155 16 159 20
rect 162 16 166 20
rect 78 11 82 15
rect 85 11 89 15
rect 92 11 96 15
rect 99 11 103 15
rect 106 11 110 15
rect 113 11 117 15
rect 120 11 124 15
rect 127 11 131 15
rect 134 11 138 15
rect 141 11 145 15
rect 148 11 152 15
rect 155 11 159 15
rect 162 11 166 15
rect 78 6 82 10
rect 85 6 89 10
rect 92 6 96 10
rect 99 6 103 10
rect 106 6 110 10
rect 113 6 117 10
rect 120 6 124 10
rect 127 6 131 10
rect 134 6 138 10
rect 141 6 145 10
rect 148 6 152 10
rect 155 6 159 10
rect 162 6 166 10
rect 9 -128 13 -124
rect 16 -128 20 -124
rect 21 -128 25 -124
rect 26 -128 30 -124
rect 31 -128 35 -124
rect 36 -128 40 -124
rect 41 -128 45 -124
rect 46 -128 50 -124
rect 51 -128 55 -124
rect 56 -128 60 -124
rect 61 -128 65 -124
rect 66 -128 70 -124
rect 73 -128 77 -124
rect 169 -128 173 -124
rect 176 -128 180 -124
rect 181 -128 185 -124
rect 186 -128 190 -124
rect 191 -128 195 -124
rect 196 -128 200 -124
rect 201 -128 205 -124
rect 206 -128 210 -124
rect 211 -128 215 -124
rect 216 -128 220 -124
rect 221 -128 225 -124
rect 226 -128 230 -124
rect 233 -128 237 -124
rect 93 -149 97 -145
rect 151 -149 155 -145
rect 93 -165 97 -161
rect 151 -165 155 -161
rect -12 -180 -8 -176
rect -7 -180 -3 -176
rect 93 -181 97 -177
rect -12 -185 -8 -181
rect -7 -185 -3 -181
rect 151 -181 155 -177
rect -12 -190 -8 -186
rect -7 -190 -3 -186
rect -12 -195 -8 -191
rect -7 -195 -3 -191
rect -12 -200 -8 -196
rect -7 -200 -3 -196
rect 93 -197 97 -193
rect -12 -205 -8 -201
rect -7 -205 -3 -201
rect -12 -210 -8 -206
rect -7 -210 -3 -206
rect -12 -215 -8 -211
rect -7 -215 -3 -211
rect -12 -220 -8 -216
rect -7 -220 -3 -216
rect -12 -225 -8 -221
rect -7 -225 -3 -221
rect -12 -230 -8 -226
rect -7 -230 -3 -226
rect -12 -235 -8 -231
rect -7 -235 -3 -231
rect -12 -240 -8 -236
rect -7 -240 -3 -236
rect 151 -197 155 -193
rect 193 -258 197 -254
rect 198 -258 202 -254
rect 203 -258 207 -254
rect 208 -258 212 -254
rect 213 -258 217 -254
rect 218 -258 222 -254
rect 223 -258 227 -254
rect 228 -258 232 -254
rect 233 -258 237 -254
rect 238 -258 242 -254
rect 243 -258 247 -254
rect 193 -263 197 -259
rect 198 -263 202 -259
rect 203 -263 207 -259
rect 208 -263 212 -259
rect 213 -263 217 -259
rect 218 -263 222 -259
rect 223 -263 227 -259
rect 228 -263 232 -259
rect 233 -263 237 -259
rect 238 -263 242 -259
rect 243 -263 247 -259
<< metal2 >>
rect 65 25 181 26
rect 65 21 78 25
rect 82 21 85 25
rect 89 21 92 25
rect 96 21 99 25
rect 103 21 106 25
rect 110 21 113 25
rect 117 21 120 25
rect 124 21 127 25
rect 131 21 134 25
rect 138 21 141 25
rect 145 21 148 25
rect 152 21 155 25
rect 159 21 162 25
rect 166 21 181 25
rect 65 20 181 21
rect 65 17 78 20
rect 75 16 78 17
rect 82 16 85 20
rect 89 16 92 20
rect 96 16 99 20
rect 103 16 106 20
rect 110 16 113 20
rect 117 16 120 20
rect 124 16 127 20
rect 131 16 134 20
rect 138 16 141 20
rect 145 16 148 20
rect 152 16 155 20
rect 159 16 162 20
rect 166 17 181 20
rect 166 16 171 17
rect 75 15 171 16
rect 75 11 78 15
rect 82 11 85 15
rect 89 11 92 15
rect 96 11 99 15
rect 103 11 106 15
rect 110 11 113 15
rect 117 11 120 15
rect 124 11 127 15
rect 131 11 134 15
rect 138 11 141 15
rect 145 11 148 15
rect 152 11 155 15
rect 159 11 162 15
rect 166 11 171 15
rect 75 10 171 11
rect 75 6 78 10
rect 82 6 85 10
rect 89 6 92 10
rect 96 6 99 10
rect 103 6 106 10
rect 110 6 113 10
rect 117 6 120 10
rect 124 6 127 10
rect 131 6 134 10
rect 138 6 141 10
rect 145 6 148 10
rect 152 6 155 10
rect 159 6 162 10
rect 166 6 171 10
rect 75 -23 171 6
rect 65 -112 181 -23
rect 13 -128 16 -124
rect 20 -128 21 -124
rect 25 -128 26 -124
rect 30 -128 31 -124
rect 35 -128 36 -124
rect 40 -128 41 -124
rect 45 -128 46 -124
rect 50 -128 51 -124
rect 55 -128 56 -124
rect 60 -128 61 -124
rect 65 -128 66 -124
rect 70 -128 73 -124
rect -24 -176 -3 -174
rect -24 -180 -22 -176
rect -18 -180 -17 -176
rect -13 -180 -12 -176
rect -8 -180 -7 -176
rect -24 -181 -3 -180
rect -24 -185 -22 -181
rect -18 -185 -17 -181
rect -13 -185 -12 -181
rect -8 -185 -7 -181
rect -24 -186 -3 -185
rect -24 -190 -22 -186
rect -18 -190 -17 -186
rect -13 -190 -12 -186
rect -8 -190 -7 -186
rect -24 -191 -3 -190
rect -24 -195 -22 -191
rect -18 -195 -17 -191
rect -13 -195 -12 -191
rect -8 -195 -7 -191
rect -24 -196 -3 -195
rect -24 -200 -22 -196
rect -18 -200 -17 -196
rect -13 -200 -12 -196
rect -8 -200 -7 -196
rect -24 -201 -3 -200
rect -24 -205 -22 -201
rect -18 -205 -17 -201
rect -13 -205 -12 -201
rect -8 -205 -7 -201
rect -24 -206 -3 -205
rect -24 -210 -22 -206
rect -18 -210 -17 -206
rect -13 -210 -12 -206
rect -8 -210 -7 -206
rect -24 -211 -3 -210
rect -24 -215 -22 -211
rect -18 -215 -17 -211
rect -13 -215 -12 -211
rect -8 -215 -7 -211
rect -24 -216 -3 -215
rect -24 -220 -22 -216
rect -18 -220 -17 -216
rect -13 -220 -12 -216
rect -8 -220 -7 -216
rect -24 -221 -3 -220
rect -24 -225 -22 -221
rect -18 -225 -17 -221
rect -13 -225 -12 -221
rect -8 -225 -7 -221
rect -24 -226 -3 -225
rect -24 -230 -22 -226
rect -18 -230 -17 -226
rect -13 -230 -12 -226
rect -8 -230 -7 -226
rect -24 -231 -3 -230
rect -24 -235 -22 -231
rect -18 -235 -17 -231
rect -13 -235 -12 -231
rect -8 -235 -7 -231
rect -24 -236 -3 -235
rect -24 -240 -22 -236
rect -18 -240 -17 -236
rect -13 -240 -12 -236
rect -8 -240 -7 -236
rect -24 -242 -3 -240
rect 9 -264 77 -128
rect 173 -128 176 -124
rect 180 -128 181 -124
rect 185 -128 186 -124
rect 190 -128 191 -124
rect 195 -128 196 -124
rect 200 -128 201 -124
rect 205 -128 206 -124
rect 210 -128 211 -124
rect 215 -128 216 -124
rect 220 -128 221 -124
rect 225 -128 226 -124
rect 230 -128 233 -124
rect 93 -161 97 -149
rect 93 -177 97 -165
rect 93 -193 97 -181
rect 151 -161 155 -149
rect 151 -177 155 -165
rect 151 -193 155 -181
rect 169 -207 237 -128
rect 169 -211 171 -207
rect 175 -211 176 -207
rect 180 -211 181 -207
rect 185 -211 186 -207
rect 190 -211 191 -207
rect 195 -211 196 -207
rect 200 -211 201 -207
rect 205 -211 206 -207
rect 210 -211 211 -207
rect 215 -211 216 -207
rect 220 -211 221 -207
rect 225 -211 226 -207
rect 230 -211 231 -207
rect 235 -211 237 -207
rect 169 -212 237 -211
rect 169 -216 171 -212
rect 175 -216 176 -212
rect 180 -216 181 -212
rect 185 -216 186 -212
rect 190 -216 191 -212
rect 195 -216 196 -212
rect 200 -216 201 -212
rect 205 -216 206 -212
rect 210 -216 211 -212
rect 215 -216 216 -212
rect 220 -216 221 -212
rect 225 -216 226 -212
rect 230 -216 231 -212
rect 235 -216 237 -212
rect 169 -219 237 -216
rect 9 -268 11 -264
rect 15 -268 16 -264
rect 20 -268 21 -264
rect 25 -268 26 -264
rect 30 -268 31 -264
rect 35 -268 36 -264
rect 40 -268 41 -264
rect 45 -268 46 -264
rect 50 -268 51 -264
rect 55 -268 56 -264
rect 60 -268 61 -264
rect 65 -268 66 -264
rect 70 -268 71 -264
rect 75 -268 77 -264
rect 9 -269 77 -268
rect 9 -273 11 -269
rect 15 -273 16 -269
rect 20 -273 21 -269
rect 25 -273 26 -269
rect 30 -273 31 -269
rect 35 -273 36 -269
rect 40 -273 41 -269
rect 45 -273 46 -269
rect 50 -273 51 -269
rect 55 -273 56 -269
rect 60 -273 61 -269
rect 65 -273 66 -269
rect 70 -273 71 -269
rect 75 -273 77 -269
rect 9 -276 77 -273
rect 197 -258 198 -254
rect 202 -258 203 -254
rect 207 -258 208 -254
rect 212 -258 213 -254
rect 217 -258 218 -254
rect 222 -258 223 -254
rect 227 -258 228 -254
rect 232 -258 233 -254
rect 237 -258 238 -254
rect 242 -258 243 -254
rect 247 -258 249 -254
rect 193 -259 249 -258
rect 197 -263 198 -259
rect 202 -263 203 -259
rect 207 -263 208 -259
rect 212 -263 213 -259
rect 217 -263 218 -259
rect 222 -263 223 -259
rect 227 -263 228 -259
rect 232 -263 233 -259
rect 237 -263 238 -259
rect 242 -263 243 -259
rect 247 -263 249 -259
rect 193 -264 249 -263
rect 197 -268 198 -264
rect 202 -268 203 -264
rect 207 -268 208 -264
rect 212 -268 213 -264
rect 217 -268 218 -264
rect 222 -268 223 -264
rect 227 -268 228 -264
rect 232 -268 233 -264
rect 237 -268 238 -264
rect 242 -268 243 -264
rect 247 -268 249 -264
rect 193 -269 249 -268
rect 197 -273 198 -269
rect 202 -273 203 -269
rect 207 -273 208 -269
rect 212 -273 213 -269
rect 217 -273 218 -269
rect 222 -273 223 -269
rect 227 -273 228 -269
rect 232 -273 233 -269
rect 237 -273 238 -269
rect 242 -273 243 -269
rect 247 -273 249 -269
rect 193 -275 249 -273
<< m3contact >>
rect -22 -180 -18 -176
rect -17 -180 -13 -176
rect -22 -185 -18 -181
rect -17 -185 -13 -181
rect -22 -190 -18 -186
rect -17 -190 -13 -186
rect -22 -195 -18 -191
rect -17 -195 -13 -191
rect -22 -200 -18 -196
rect -17 -200 -13 -196
rect -22 -205 -18 -201
rect -17 -205 -13 -201
rect -22 -210 -18 -206
rect -17 -210 -13 -206
rect -22 -215 -18 -211
rect -17 -215 -13 -211
rect -22 -220 -18 -216
rect -17 -220 -13 -216
rect -22 -225 -18 -221
rect -17 -225 -13 -221
rect -22 -230 -18 -226
rect -17 -230 -13 -226
rect -22 -235 -18 -231
rect -17 -235 -13 -231
rect -22 -240 -18 -236
rect -17 -240 -13 -236
rect 171 -211 175 -207
rect 176 -211 180 -207
rect 181 -211 185 -207
rect 186 -211 190 -207
rect 191 -211 195 -207
rect 196 -211 200 -207
rect 201 -211 205 -207
rect 206 -211 210 -207
rect 211 -211 215 -207
rect 216 -211 220 -207
rect 221 -211 225 -207
rect 226 -211 230 -207
rect 231 -211 235 -207
rect 171 -216 175 -212
rect 176 -216 180 -212
rect 181 -216 185 -212
rect 186 -216 190 -212
rect 191 -216 195 -212
rect 196 -216 200 -212
rect 201 -216 205 -212
rect 206 -216 210 -212
rect 211 -216 215 -212
rect 216 -216 220 -212
rect 221 -216 225 -212
rect 226 -216 230 -212
rect 231 -216 235 -212
rect 11 -268 15 -264
rect 16 -268 20 -264
rect 21 -268 25 -264
rect 26 -268 30 -264
rect 31 -268 35 -264
rect 36 -268 40 -264
rect 41 -268 45 -264
rect 46 -268 50 -264
rect 51 -268 55 -264
rect 56 -268 60 -264
rect 61 -268 65 -264
rect 66 -268 70 -264
rect 71 -268 75 -264
rect 11 -273 15 -269
rect 16 -273 20 -269
rect 21 -273 25 -269
rect 26 -273 30 -269
rect 31 -273 35 -269
rect 36 -273 40 -269
rect 41 -273 45 -269
rect 46 -273 50 -269
rect 51 -273 55 -269
rect 56 -273 60 -269
rect 61 -273 65 -269
rect 66 -273 70 -269
rect 71 -273 75 -269
rect 193 -268 197 -264
rect 198 -268 202 -264
rect 203 -268 207 -264
rect 208 -268 212 -264
rect 213 -268 217 -264
rect 218 -268 222 -264
rect 223 -268 227 -264
rect 228 -268 232 -264
rect 233 -268 237 -264
rect 238 -268 242 -264
rect 243 -268 247 -264
rect 193 -273 197 -269
rect 198 -273 202 -269
rect 203 -273 207 -269
rect 208 -273 212 -269
rect 213 -273 217 -269
rect 218 -273 222 -269
rect 223 -273 227 -269
rect 228 -273 232 -269
rect 233 -273 237 -269
rect 238 -273 242 -269
rect 243 -273 247 -269
<< metal3 >>
rect -24 -176 -12 -174
rect -24 -180 -22 -176
rect -18 -180 -17 -176
rect -13 -180 -12 -176
rect -24 -181 -12 -180
rect -24 -185 -22 -181
rect -18 -185 -17 -181
rect -13 -185 -12 -181
rect -24 -186 -12 -185
rect -24 -190 -22 -186
rect -18 -190 -17 -186
rect -13 -190 -12 -186
rect -24 -191 -12 -190
rect -24 -195 -22 -191
rect -18 -195 -17 -191
rect -13 -195 -12 -191
rect -24 -196 -12 -195
rect -24 -200 -22 -196
rect -18 -200 -17 -196
rect -13 -200 -12 -196
rect -24 -201 -12 -200
rect -24 -205 -22 -201
rect -18 -205 -17 -201
rect -13 -205 -12 -201
rect -24 -206 -12 -205
rect -24 -210 -22 -206
rect -18 -210 -17 -206
rect -13 -210 -12 -206
rect -24 -211 -12 -210
rect -24 -215 -22 -211
rect -18 -215 -17 -211
rect -13 -215 -12 -211
rect -24 -216 -12 -215
rect -24 -220 -22 -216
rect -18 -220 -17 -216
rect -13 -220 -12 -216
rect 169 -207 237 -206
rect 169 -211 171 -207
rect 175 -211 176 -207
rect 180 -211 181 -207
rect 185 -211 186 -207
rect 190 -211 191 -207
rect 195 -211 196 -207
rect 200 -211 201 -207
rect 205 -211 206 -207
rect 210 -211 211 -207
rect 215 -211 216 -207
rect 220 -211 221 -207
rect 225 -211 226 -207
rect 230 -211 231 -207
rect 235 -211 237 -207
rect 169 -212 237 -211
rect 169 -216 171 -212
rect 175 -216 176 -212
rect 180 -216 181 -212
rect 185 -216 186 -212
rect 190 -216 191 -212
rect 195 -216 196 -212
rect 200 -216 201 -212
rect 205 -216 206 -212
rect 210 -216 211 -212
rect 215 -216 216 -212
rect 220 -216 221 -212
rect 225 -216 226 -212
rect 230 -216 231 -212
rect 235 -216 237 -212
rect 169 -219 237 -216
rect -24 -221 -12 -220
rect -24 -225 -22 -221
rect -18 -225 -17 -221
rect -13 -225 -12 -221
rect -24 -226 -12 -225
rect -24 -230 -22 -226
rect -18 -230 -17 -226
rect -13 -230 -12 -226
rect -24 -231 -12 -230
rect -24 -235 -22 -231
rect -18 -235 -17 -231
rect -13 -235 -12 -231
rect -24 -236 -12 -235
rect -24 -240 -22 -236
rect -18 -240 -17 -236
rect -13 -240 -12 -236
rect -24 -243 -12 -240
rect 9 -264 77 -263
rect 9 -268 11 -264
rect 15 -268 16 -264
rect 20 -268 21 -264
rect 25 -268 26 -264
rect 30 -268 31 -264
rect 35 -268 36 -264
rect 40 -268 41 -264
rect 45 -268 46 -264
rect 50 -268 51 -264
rect 55 -268 56 -264
rect 60 -268 61 -264
rect 65 -268 66 -264
rect 70 -268 71 -264
rect 75 -268 77 -264
rect 9 -269 77 -268
rect 9 -273 11 -269
rect 15 -273 16 -269
rect 20 -273 21 -269
rect 25 -273 26 -269
rect 30 -273 31 -269
rect 35 -273 36 -269
rect 40 -273 41 -269
rect 45 -273 46 -269
rect 50 -273 51 -269
rect 55 -273 56 -269
rect 60 -273 61 -269
rect 65 -273 66 -269
rect 70 -273 71 -269
rect 75 -273 77 -269
rect 9 -276 77 -273
rect 192 -264 249 -262
rect 192 -268 193 -264
rect 197 -268 198 -264
rect 202 -268 203 -264
rect 207 -268 208 -264
rect 212 -268 213 -264
rect 217 -268 218 -264
rect 222 -268 223 -264
rect 227 -268 228 -264
rect 232 -268 233 -264
rect 237 -268 238 -264
rect 242 -268 243 -264
rect 247 -268 249 -264
rect 192 -269 249 -268
rect 192 -273 193 -269
rect 197 -273 198 -269
rect 202 -273 203 -269
rect 207 -273 208 -269
rect 212 -273 213 -269
rect 217 -273 218 -269
rect 222 -273 223 -269
rect 227 -273 228 -269
rect 232 -273 233 -269
rect 237 -273 238 -269
rect 242 -273 243 -269
rect 247 -273 249 -269
rect 192 -275 249 -273
use barepad  b
timestamp 1006127261
transform 1 0 -23 0 1 -697
box 16 702 276 1014
use ndiode  nd
timestamp 1037203521
transform 1 0 9 0 1 -125
box -14 -13 82 128
use pdiode  pd
timestamp 1037203492
transform 1 0 148 0 1 -129
box 7 -9 103 132
use barering  br
timestamp 1006127261
transform 1 0 -34 0 1 -343
box 2 -23 311 176
<< labels >>
rlabel metal3 -17 -237 -17 -237 1 Vdd!
rlabel metal1 123 -122 123 -122 1 RawIn
rlabel metal1 122 -200 122 -200 1 in
rlabel metal1 116 -155 116 -155 1 _RawIn
<< end >>
