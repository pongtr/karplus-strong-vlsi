magic
tech scmos
timestamp 1512712928
<< nwell >>
rect -27 -9 2 9
<< pwell >>
rect -32 -27 -3 -9
<< ntransistor >>
rect -16 -18 -14 -15
<< ptransistor >>
rect -16 -3 -14 3
<< ndiffusion >>
rect -17 -18 -16 -15
rect -14 -18 -13 -15
<< pdiffusion >>
rect -17 -3 -16 3
rect -14 1 -9 3
rect -14 -3 -13 1
<< ndcontact >>
rect -21 -19 -17 -15
rect -13 -19 -9 -15
<< pdcontact >>
rect -21 -3 -17 3
rect -13 -3 -9 1
<< psubstratepcontact >>
rect -29 -23 -25 -19
<< nsubstratencontact >>
rect -5 1 -1 5
<< polysilicon >>
rect -16 3 -14 5
rect -16 -15 -14 -3
rect -16 -20 -14 -18
<< polycontact >>
rect -20 -11 -16 -7
<< metal1 >>
rect -13 -7 -9 -3
rect -32 -11 -20 -7
rect -13 -11 3 -7
rect -13 -15 -9 -11
<< m2contact >>
rect -25 -3 -21 1
rect -5 -3 -1 1
rect -29 -19 -25 -15
rect -21 -23 -17 -19
<< metal2 >>
rect -29 -15 -25 1
rect -5 -19 -1 -3
rect -17 -23 -1 -19
<< labels >>
rlabel m2contact -27 -17 -27 -17 3 Vdd
<< end >>
